magic
tech scmos
timestamp 1681685098
<< metal1 >>
rect 14 2007 2204 2027
rect 38 1983 2180 2003
rect 38 1967 2180 1973
rect 508 1943 517 1946
rect 1098 1943 1108 1946
rect 228 1933 269 1936
rect 274 1926 277 1935
rect 500 1933 541 1936
rect 562 1926 565 1935
rect 618 1926 621 1935
rect 692 1933 717 1936
rect 874 1933 884 1936
rect 1012 1933 1044 1936
rect 1092 1933 1116 1936
rect 1138 1926 1141 1935
rect 1188 1933 1196 1936
rect 1338 1933 1348 1936
rect 1378 1926 1381 1935
rect 1428 1933 1437 1936
rect 1450 1933 1460 1936
rect 1660 1933 1676 1936
rect 1826 1933 1860 1936
rect 1900 1933 1917 1936
rect 2018 1926 2021 1935
rect 162 1923 172 1926
rect 242 1923 277 1926
rect 394 1923 412 1926
rect 450 1923 484 1926
rect 562 1923 588 1926
rect 618 1923 676 1926
rect 706 1923 724 1926
rect 836 1923 892 1926
rect 1018 1923 1060 1926
rect 1132 1923 1141 1926
rect 1204 1923 1220 1926
rect 1364 1923 1381 1926
rect 1476 1923 1500 1926
rect 1532 1923 1557 1926
rect 1708 1923 1725 1926
rect 1762 1923 1788 1926
rect 1882 1923 1892 1926
rect 1956 1923 1981 1926
rect 2012 1923 2021 1926
rect 2028 1923 2044 1926
rect 538 1913 548 1916
rect 1434 1913 1460 1916
rect 1546 1913 1564 1916
rect 1578 1913 1588 1916
rect 2060 1913 2069 1916
rect 14 1867 2204 1873
rect 308 1823 333 1826
rect 914 1823 932 1826
rect 1146 1823 1156 1826
rect 1370 1823 1396 1826
rect 1754 1816 1757 1825
rect 1946 1823 1964 1826
rect 188 1813 197 1816
rect 108 1803 125 1806
rect 162 1803 172 1806
rect 202 1803 205 1814
rect 218 1813 285 1816
rect 500 1813 525 1816
rect 556 1813 565 1816
rect 580 1813 644 1816
rect 676 1813 701 1816
rect 796 1813 821 1816
rect 908 1813 925 1816
rect 948 1813 965 1816
rect 1004 1813 1013 1816
rect 1164 1813 1181 1816
rect 1194 1813 1204 1816
rect 1404 1813 1437 1816
rect 236 1803 245 1806
rect 282 1803 285 1813
rect 386 1803 396 1806
rect 652 1803 661 1806
rect 682 1803 780 1806
rect 386 1795 389 1803
rect 658 1795 661 1803
rect 1578 1796 1581 1814
rect 1674 1813 1740 1816
rect 1754 1813 1772 1816
rect 1876 1813 1885 1816
rect 1938 1813 1972 1816
rect 2020 1813 2037 1816
rect 2052 1813 2069 1816
rect 1642 1803 1652 1806
rect 1714 1803 1732 1806
rect 2036 1803 2045 1806
rect 796 1793 884 1796
rect 1578 1793 1644 1796
rect 38 1767 2180 1773
rect 122 1743 188 1746
rect 482 1743 548 1746
rect 682 1743 708 1746
rect 1148 1743 1181 1746
rect 82 1733 92 1736
rect 154 1723 157 1743
rect 682 1736 685 1743
rect 218 1726 221 1735
rect 212 1723 221 1726
rect 282 1725 285 1736
rect 388 1733 397 1736
rect 426 1733 436 1736
rect 668 1733 685 1736
rect 738 1726 741 1735
rect 1010 1733 1020 1736
rect 1140 1733 1157 1736
rect 346 1723 372 1726
rect 452 1723 468 1726
rect 572 1723 621 1726
rect 732 1723 741 1726
rect 812 1723 844 1726
rect 898 1723 916 1726
rect 1036 1723 1125 1726
rect 1234 1716 1237 1736
rect 1242 1733 1292 1736
rect 1612 1733 1620 1736
rect 1762 1726 1765 1735
rect 1850 1733 1876 1736
rect 1970 1733 1980 1736
rect 2028 1733 2044 1736
rect 1282 1723 1300 1726
rect 1444 1723 1453 1726
rect 1540 1723 1557 1726
rect 1708 1723 1765 1726
rect 1892 1723 1909 1726
rect 1930 1723 1956 1726
rect 1978 1723 1996 1726
rect 116 1713 133 1716
rect 276 1713 285 1716
rect 300 1713 325 1716
rect 578 1713 628 1716
rect 924 1713 965 1716
rect 1002 1713 1020 1716
rect 1220 1713 1237 1716
rect 1316 1713 1389 1716
rect 1794 1713 1876 1716
rect 274 1703 292 1706
rect 1154 1703 1212 1706
rect 14 1667 2204 1673
rect 330 1623 356 1626
rect 658 1623 684 1626
rect 962 1623 996 1626
rect 1410 1623 1444 1626
rect 1620 1623 1629 1626
rect 1626 1616 1629 1623
rect 130 1613 140 1616
rect 146 1613 172 1616
rect 266 1613 292 1616
rect 364 1613 381 1616
rect 420 1613 429 1616
rect 482 1613 492 1616
rect 650 1613 692 1616
rect 698 1613 724 1616
rect 796 1613 805 1616
rect 1010 1613 1036 1616
rect 1164 1613 1189 1616
rect 1226 1613 1236 1616
rect 1314 1613 1332 1616
rect 1386 1613 1396 1616
rect 1452 1613 1469 1616
rect 1532 1613 1541 1616
rect 556 1603 581 1606
rect 698 1605 701 1613
rect 882 1603 892 1606
rect 940 1603 949 1606
rect 1010 1605 1013 1613
rect 1068 1603 1077 1606
rect 1258 1603 1268 1606
rect 1314 1605 1317 1613
rect 1378 1603 1388 1606
rect 1594 1605 1597 1616
rect 1626 1613 1644 1616
rect 1724 1613 1756 1616
rect 1844 1613 1853 1616
rect 1906 1613 1916 1616
rect 2004 1613 2021 1616
rect 2060 1613 2069 1616
rect 1738 1603 1748 1606
rect 506 1593 548 1596
rect 882 1595 885 1603
rect 1258 1595 1261 1603
rect 2066 1596 2069 1613
rect 2066 1593 2100 1596
rect 38 1567 2180 1573
rect 556 1543 565 1546
rect 1746 1543 1788 1546
rect 1890 1543 1900 1546
rect 1890 1536 1893 1543
rect 372 1533 397 1536
rect 436 1533 452 1536
rect 698 1533 708 1536
rect 732 1533 757 1536
rect 1130 1533 1140 1536
rect 1186 1533 1228 1536
rect 394 1526 397 1533
rect 1250 1526 1253 1535
rect 1340 1533 1373 1536
rect 1378 1533 1396 1536
rect 1450 1533 1469 1536
rect 1500 1533 1509 1536
rect 108 1523 117 1526
rect 196 1523 253 1526
rect 276 1523 285 1526
rect 346 1523 356 1526
rect 394 1523 420 1526
rect 484 1523 501 1526
rect 506 1523 532 1526
rect 684 1523 693 1526
rect 698 1523 716 1526
rect 914 1523 972 1526
rect 1026 1523 1052 1526
rect 1148 1523 1157 1526
rect 1250 1523 1261 1526
rect 1322 1523 1332 1526
rect 1362 1523 1469 1526
rect 1506 1523 1580 1526
rect 1698 1523 1708 1526
rect 1818 1523 1821 1535
rect 1868 1533 1893 1536
rect 1898 1533 1908 1536
rect 2060 1533 2084 1536
rect 2132 1533 2141 1536
rect 1924 1523 1957 1526
rect 1994 1523 2004 1526
rect 2018 1523 2036 1526
rect 2058 1523 2100 1526
rect 1258 1516 1261 1523
rect 218 1513 260 1516
rect 732 1513 829 1516
rect 834 1513 884 1516
rect 908 1513 933 1516
rect 1218 1513 1228 1516
rect 1258 1513 1292 1516
rect 1938 1513 1964 1516
rect 2018 1515 2021 1523
rect 14 1467 2204 1473
rect 1460 1433 1469 1436
rect 428 1423 453 1426
rect 972 1423 1013 1426
rect 1210 1423 1228 1426
rect 1282 1423 1332 1426
rect 1394 1423 1412 1426
rect 1442 1423 1452 1426
rect 1700 1423 1709 1426
rect 1714 1423 1788 1426
rect 2060 1423 2069 1426
rect 1442 1416 1445 1423
rect 108 1413 133 1416
rect 164 1413 173 1416
rect 282 1413 292 1416
rect 258 1403 284 1406
rect 338 1403 356 1406
rect 402 1405 405 1416
rect 516 1413 541 1416
rect 538 1405 541 1413
rect 626 1413 700 1416
rect 884 1413 909 1416
rect 986 1413 1020 1416
rect 1066 1413 1148 1416
rect 1244 1413 1253 1416
rect 1340 1413 1413 1416
rect 1434 1413 1445 1416
rect 626 1403 629 1413
rect 994 1403 1012 1406
rect 1026 1403 1036 1406
rect 1090 1403 1140 1406
rect 1164 1403 1181 1406
rect 1218 1403 1228 1406
rect 1252 1403 1269 1406
rect 1434 1405 1437 1413
rect 1466 1403 1469 1414
rect 1530 1413 1556 1416
rect 1668 1413 1684 1416
rect 1650 1403 1660 1406
rect 1794 1403 1797 1414
rect 1882 1413 1900 1416
rect 1956 1413 1981 1416
rect 2012 1413 2021 1416
rect 2028 1413 2044 1416
rect 1842 1403 1908 1406
rect 2018 1405 2021 1413
rect 1844 1393 1901 1396
rect 38 1367 2180 1373
rect 300 1343 317 1346
rect 738 1343 748 1346
rect 738 1336 741 1343
rect 1042 1336 1045 1345
rect 1786 1343 1796 1346
rect 244 1335 269 1336
rect 242 1333 269 1335
rect 292 1333 325 1336
rect 108 1323 117 1326
rect 242 1323 245 1333
rect 530 1326 533 1335
rect 716 1333 741 1336
rect 778 1326 781 1335
rect 914 1333 940 1336
rect 954 1326 957 1336
rect 1036 1333 1045 1336
rect 1052 1333 1061 1336
rect 1138 1326 1141 1335
rect 1258 1333 1268 1336
rect 1290 1335 1316 1336
rect 1290 1333 1317 1335
rect 1506 1333 1524 1336
rect 1588 1333 1605 1336
rect 1610 1333 1636 1336
rect 1314 1326 1317 1333
rect 1690 1326 1693 1335
rect 1706 1333 1732 1336
rect 1786 1333 1804 1336
rect 274 1323 284 1326
rect 332 1323 357 1326
rect 468 1323 493 1326
rect 524 1323 533 1326
rect 540 1323 549 1326
rect 658 1323 676 1326
rect 772 1323 781 1326
rect 812 1323 837 1326
rect 954 1323 1028 1326
rect 1060 1323 1069 1326
rect 1138 1323 1148 1326
rect 1178 1323 1204 1326
rect 1314 1323 1333 1326
rect 1498 1323 1548 1326
rect 1562 1323 1580 1326
rect 1668 1323 1693 1326
rect 1834 1326 1837 1335
rect 2018 1326 2021 1335
rect 2034 1333 2052 1336
rect 1834 1323 1852 1326
rect 1882 1323 1908 1326
rect 1996 1323 2021 1326
rect 2068 1323 2141 1326
rect 354 1316 357 1323
rect 354 1313 372 1316
rect 636 1313 645 1316
rect 834 1313 884 1316
rect 908 1313 917 1316
rect 346 1303 388 1306
rect 1066 1303 1069 1323
rect 1074 1313 1124 1316
rect 1562 1315 1565 1323
rect 1708 1313 1725 1316
rect 14 1267 2204 1273
rect 234 1216 237 1225
rect 708 1223 733 1226
rect 964 1223 1021 1226
rect 146 1213 172 1216
rect 220 1213 237 1216
rect 252 1213 269 1216
rect 314 1213 332 1216
rect 474 1213 484 1216
rect 530 1213 540 1216
rect 642 1213 692 1216
rect 786 1213 796 1216
rect 850 1213 885 1216
rect 962 1213 1036 1216
rect 1164 1213 1181 1216
rect 850 1206 853 1213
rect 1394 1206 1397 1216
rect 1548 1213 1565 1216
rect 1676 1213 1709 1216
rect 1722 1213 1732 1216
rect 1762 1207 1765 1216
rect 1772 1213 1813 1216
rect 1834 1213 1845 1216
rect 2028 1213 2053 1216
rect 1834 1207 1837 1213
rect 108 1203 156 1206
rect 316 1203 324 1206
rect 610 1203 620 1206
rect 674 1203 684 1206
rect 788 1203 797 1206
rect 812 1203 853 1206
rect 858 1203 868 1206
rect 914 1203 940 1206
rect 1044 1203 1053 1206
rect 1082 1203 1140 1206
rect 1170 1203 1180 1206
rect 1292 1203 1325 1206
rect 1388 1203 1397 1206
rect 1610 1203 1660 1206
rect 586 1193 612 1196
rect 1050 1195 1053 1203
rect 1754 1195 1757 1206
rect 1802 1203 1812 1206
rect 1954 1203 1972 1206
rect 1946 1193 1964 1196
rect 38 1167 2180 1173
rect 1588 1143 1597 1146
rect 82 1133 92 1136
rect 130 1123 156 1126
rect 162 1123 196 1126
rect 338 1123 341 1134
rect 388 1133 405 1136
rect 548 1133 581 1136
rect 636 1133 661 1136
rect 804 1133 844 1136
rect 354 1123 364 1126
rect 530 1123 540 1126
rect 546 1123 612 1126
rect 700 1123 709 1126
rect 796 1123 805 1126
rect 810 1123 852 1126
rect 890 1123 1020 1126
rect 1026 1123 1029 1134
rect 1106 1133 1116 1136
rect 1164 1133 1173 1136
rect 1330 1133 1356 1136
rect 1466 1133 1476 1136
rect 1562 1133 1580 1136
rect 1660 1133 1717 1136
rect 1746 1133 1756 1136
rect 1876 1133 1885 1136
rect 1562 1126 1565 1133
rect 1052 1123 1077 1126
rect 1130 1123 1140 1126
rect 1204 1123 1237 1126
rect 1260 1123 1293 1126
rect 1324 1123 1357 1126
rect 1380 1123 1469 1126
rect 1516 1123 1565 1126
rect 1586 1123 1685 1126
rect 1826 1123 1836 1126
rect 1874 1123 1916 1126
rect 2026 1123 2036 1126
rect 130 1116 133 1123
rect 116 1113 133 1116
rect 138 1113 148 1116
rect 1876 1113 1909 1116
rect 2044 1113 2061 1116
rect 14 1067 2204 1073
rect 1732 1033 1749 1036
rect 484 1023 493 1026
rect 1674 1023 1724 1026
rect 1748 1023 1796 1026
rect 1810 1023 1820 1026
rect 186 1013 212 1016
rect 452 1013 468 1016
rect 482 1013 516 1016
rect 772 1013 789 1016
rect 828 1013 869 1016
rect 874 1013 900 1016
rect 1146 1013 1180 1016
rect 1316 1013 1349 1016
rect 1538 1013 1548 1016
rect 1554 1013 1564 1016
rect 1668 1013 1717 1016
rect 1786 1013 1804 1016
rect 1554 1007 1557 1013
rect 2050 1006 2053 1014
rect 242 1003 260 1006
rect 498 1003 524 1006
rect 602 1003 620 1006
rect 882 1003 892 1006
rect 1202 1003 1212 1006
rect 1324 1003 1341 1006
rect 1466 1003 1492 1006
rect 2034 1003 2044 1006
rect 2050 1003 2117 1006
rect 554 993 612 996
rect 38 967 2180 973
rect 266 933 292 936
rect 322 933 364 936
rect 404 933 461 936
rect 602 933 612 936
rect 700 933 733 936
rect 834 933 868 936
rect 1052 933 1061 936
rect 1210 933 1260 936
rect 1460 933 1517 936
rect 1684 933 1757 936
rect 1836 933 1845 936
rect 1972 933 1981 936
rect 148 923 157 926
rect 372 923 381 926
rect 418 923 460 926
rect 522 923 548 926
rect 636 923 669 926
rect 804 923 925 926
rect 978 923 1036 926
rect 1058 923 1164 926
rect 1196 923 1261 926
rect 1306 923 1309 933
rect 1340 923 1349 926
rect 1490 923 1493 933
rect 1842 926 1845 933
rect 1514 923 1540 926
rect 1818 923 1828 926
rect 1842 923 1852 926
rect 2108 923 2117 926
rect 2132 923 2149 926
rect 922 916 925 923
rect 922 913 956 916
rect 1052 913 1069 916
rect 1786 913 1804 916
rect 2114 915 2117 923
rect 14 867 2204 873
rect 666 833 676 836
rect 642 823 660 826
rect 684 823 741 826
rect 1588 823 1645 826
rect 1820 823 1828 826
rect 2044 823 2069 826
rect 116 813 157 816
rect 180 813 189 816
rect 298 813 317 816
rect 322 813 380 816
rect 564 813 581 816
rect 602 813 612 816
rect 690 813 756 816
rect 786 813 836 816
rect 996 813 1005 816
rect 1034 813 1084 816
rect 1090 813 1100 816
rect 1172 813 1197 816
rect 154 807 157 813
rect 314 807 317 813
rect 1258 807 1261 816
rect 1354 813 1373 816
rect 1514 813 1572 816
rect 1370 807 1373 813
rect 1586 807 1589 816
rect 1668 813 1716 816
rect 1738 813 1812 816
rect 1818 813 1836 816
rect 1924 813 1949 816
rect 1980 813 1997 816
rect 2012 813 2021 816
rect 2058 813 2116 816
rect 82 803 92 806
rect 316 803 373 806
rect 404 803 437 806
rect 442 803 460 806
rect 508 803 524 806
rect 556 803 613 806
rect 620 803 653 806
rect 780 803 797 806
rect 826 803 844 806
rect 1124 803 1133 806
rect 1154 803 1164 806
rect 1314 803 1324 806
rect 1538 803 1564 806
rect 1642 803 1652 806
rect 1732 803 1749 806
rect 1786 803 1804 806
rect 1986 803 2004 806
rect 2010 803 2020 806
rect 2044 803 2053 806
rect 38 767 2180 773
rect 650 743 676 746
rect 1218 743 1229 746
rect 1738 743 1796 746
rect 1226 736 1229 743
rect 180 733 188 736
rect 562 733 580 736
rect 642 733 684 736
rect 868 733 973 736
rect 988 733 1013 736
rect 1098 733 1140 736
rect 1164 733 1221 736
rect 1226 733 1236 736
rect 1010 726 1013 733
rect 108 723 149 726
rect 212 723 261 726
rect 420 723 436 726
rect 692 723 749 726
rect 962 723 972 726
rect 996 723 1005 726
rect 1010 723 1084 726
rect 1156 723 1181 726
rect 1338 723 1341 734
rect 1442 733 1468 736
rect 1530 733 1588 736
rect 1618 733 1628 736
rect 1666 733 1692 736
rect 1804 733 1813 736
rect 1850 733 1876 736
rect 1362 723 1428 726
rect 1484 723 1493 726
rect 1604 723 1629 726
rect 1636 723 1685 726
rect 1700 723 1709 726
rect 1812 723 1820 726
rect 1844 723 1861 726
rect 1866 723 1884 726
rect 1954 723 1980 726
rect 2108 723 2117 726
rect 1364 713 1397 716
rect 1402 713 1420 716
rect 1434 713 1468 716
rect 1514 713 1524 716
rect 1402 706 1405 713
rect 1370 703 1405 706
rect 14 667 2204 673
rect 788 623 813 626
rect 1348 623 1373 626
rect 1644 623 1677 626
rect 1370 616 1373 623
rect 82 613 92 616
rect 186 607 189 616
rect 268 613 277 616
rect 306 613 325 616
rect 412 613 429 616
rect 780 613 861 616
rect 890 613 948 616
rect 972 613 989 616
rect 1068 613 1172 616
rect 1218 613 1245 616
rect 1340 613 1365 616
rect 1370 613 1404 616
rect 1636 613 1765 616
rect 274 607 277 613
rect 322 607 325 613
rect 1242 607 1245 613
rect 2122 607 2125 616
rect 2132 613 2149 616
rect 330 603 364 606
rect 404 603 469 606
rect 500 603 533 606
rect 620 603 637 606
rect 762 603 772 606
rect 884 603 949 606
rect 970 603 1052 606
rect 1076 603 1133 606
rect 1138 603 1164 606
rect 1346 603 1396 606
rect 1514 603 1628 606
rect 530 593 540 596
rect 946 595 949 603
rect 38 567 2180 573
rect 220 533 229 536
rect 388 533 397 536
rect 420 533 445 536
rect 564 533 580 536
rect 914 533 924 536
rect 948 533 957 536
rect 1188 533 1252 536
rect 1266 533 1308 536
rect 1554 533 1564 536
rect 1626 533 1660 536
rect 1676 533 1693 536
rect 1828 533 1861 536
rect 1892 533 1917 536
rect 2052 533 2061 536
rect 2108 533 2117 536
rect 682 526 685 533
rect 890 526 893 533
rect 386 523 396 526
rect 626 523 685 526
rect 724 523 732 526
rect 890 523 932 526
rect 994 523 1020 526
rect 1058 523 1156 526
rect 1162 523 1172 526
rect 1250 523 1260 526
rect 1266 523 1269 533
rect 1418 523 1421 533
rect 1530 526 1533 533
rect 1922 526 1925 533
rect 1468 523 1493 526
rect 1524 523 1533 526
rect 1540 523 1572 526
rect 1594 523 1652 526
rect 1708 523 1781 526
rect 1786 523 1820 526
rect 1884 523 1901 526
rect 1906 523 1925 526
rect 1946 526 1949 533
rect 2074 526 2077 533
rect 1946 523 1957 526
rect 1970 523 2012 526
rect 2050 523 2077 526
rect 826 513 876 516
rect 1588 513 1613 516
rect 1826 513 1876 516
rect 1978 513 2004 516
rect 2052 513 2069 516
rect 14 467 2204 473
rect 876 423 909 426
rect 1452 423 1477 426
rect 1700 423 1709 426
rect 1714 423 1740 426
rect 1786 423 1804 426
rect 1882 416 1885 425
rect 2066 423 2092 426
rect 108 413 149 416
rect 212 413 261 416
rect 388 413 404 416
rect 508 413 524 416
rect 626 413 652 416
rect 844 413 860 416
rect 930 413 948 416
rect 1018 413 1036 416
rect 1146 413 1156 416
rect 1170 413 1180 416
rect 1250 413 1260 416
rect 1396 413 1436 416
rect 1490 413 1500 416
rect 1532 413 1564 416
rect 1692 413 1741 416
rect 1748 413 1789 416
rect 1868 413 1885 416
rect 138 403 156 406
rect 362 403 372 406
rect 482 403 492 406
rect 596 403 621 406
rect 730 403 836 406
rect 956 403 1020 406
rect 1114 403 1148 406
rect 1188 403 1252 406
rect 1404 403 1421 406
rect 1466 403 1508 406
rect 1530 403 1540 406
rect 1602 403 1628 406
rect 1786 403 1789 413
rect 1794 403 1804 406
rect 1828 403 1837 406
rect 1842 403 1860 406
rect 1218 393 1221 403
rect 38 367 2180 373
rect 772 343 813 346
rect 196 333 213 336
rect 244 333 261 336
rect 378 333 388 336
rect 404 333 413 336
rect 524 333 557 336
rect 562 333 572 336
rect 618 326 621 334
rect 668 333 685 336
rect 764 333 821 336
rect 682 326 685 333
rect 826 326 829 334
rect 82 323 100 326
rect 202 323 220 326
rect 250 323 380 326
rect 412 323 429 326
rect 442 323 500 326
rect 538 323 588 326
rect 618 323 652 326
rect 682 323 748 326
rect 810 323 829 326
rect 874 326 877 334
rect 972 333 1029 336
rect 1226 333 1300 336
rect 1316 333 1357 336
rect 1524 333 1565 336
rect 1596 333 1669 336
rect 1562 326 1565 333
rect 874 323 956 326
rect 1060 323 1085 326
rect 1164 323 1173 326
rect 1282 323 1292 326
rect 1420 323 1445 326
rect 1482 323 1500 326
rect 1562 323 1572 326
rect 1684 323 1773 326
rect 1780 323 1789 326
rect 1882 323 1900 326
rect 2020 323 2045 326
rect 2124 323 2133 326
rect 1692 313 1709 316
rect 14 267 2204 273
rect 1692 223 1701 226
rect 1946 216 1949 225
rect 2074 216 2077 225
rect 202 213 236 216
rect 386 205 389 216
rect 474 213 532 216
rect 586 213 620 216
rect 658 213 708 216
rect 788 213 821 216
rect 978 206 981 216
rect 986 213 1020 216
rect 1082 213 1092 216
rect 1122 213 1164 216
rect 1234 213 1252 216
rect 1282 213 1308 216
rect 420 203 501 206
rect 570 203 628 206
rect 732 203 764 206
rect 842 203 900 206
rect 946 203 996 206
rect 1188 203 1245 206
rect 1330 205 1333 216
rect 1338 213 1372 216
rect 1452 213 1485 216
rect 1684 213 1709 216
rect 1716 213 1733 216
rect 1796 213 1813 216
rect 1850 213 1932 216
rect 1946 213 1964 216
rect 1978 213 2060 216
rect 2074 213 2092 216
rect 1396 203 1428 206
rect 1482 205 1485 213
rect 1618 203 1676 206
rect 1778 203 1788 206
rect 1858 203 1924 206
rect 1970 203 2052 206
rect 38 167 2180 173
rect 122 133 132 136
rect 210 133 228 136
rect 308 133 333 136
rect 474 133 484 136
rect 564 133 573 136
rect 578 133 596 136
rect 708 133 740 136
rect 956 133 1005 136
rect 1036 133 1053 136
rect 1178 133 1204 136
rect 1378 133 1404 136
rect 1482 133 1500 136
rect 1548 133 1557 136
rect 1562 133 1572 136
rect 1666 133 1684 136
rect 162 123 180 126
rect 354 123 357 133
rect 1378 126 1381 133
rect 402 123 444 126
rect 586 123 620 126
rect 674 123 684 126
rect 764 123 797 126
rect 898 123 932 126
rect 962 123 1012 126
rect 1042 123 1060 126
rect 1090 123 1116 126
rect 1364 123 1381 126
rect 1434 123 1452 126
rect 1524 123 1549 126
rect 1554 123 1557 133
rect 1762 126 1765 133
rect 1692 123 1765 126
rect 1946 123 1964 126
rect 2068 123 2077 126
rect 14 67 2204 73
rect 38 37 2180 57
rect 14 13 2204 33
<< metal2 >>
rect 14 13 34 2027
rect 38 37 58 2003
rect 114 1923 117 1946
rect 226 1943 237 1946
rect 82 1733 85 1786
rect 98 1723 101 1816
rect 122 1743 125 1806
rect 162 1803 165 1926
rect 194 1923 197 1936
rect 234 1926 237 1943
rect 266 1933 269 1946
rect 322 1933 325 1946
rect 210 1836 213 1926
rect 234 1923 245 1926
rect 234 1856 237 1923
rect 234 1853 245 1856
rect 210 1833 229 1836
rect 170 1823 181 1826
rect 194 1823 221 1826
rect 194 1813 197 1823
rect 218 1813 221 1823
rect 194 1783 197 1806
rect 202 1776 205 1806
rect 186 1773 205 1776
rect 186 1743 189 1773
rect 114 1706 117 1736
rect 106 1703 117 1706
rect 106 1596 109 1703
rect 130 1613 133 1716
rect 146 1623 149 1636
rect 146 1606 149 1616
rect 130 1603 149 1606
rect 106 1593 117 1596
rect 82 1333 85 1546
rect 114 1523 117 1593
rect 154 1576 157 1726
rect 194 1706 197 1766
rect 210 1713 213 1806
rect 218 1783 221 1796
rect 226 1763 229 1833
rect 242 1803 245 1853
rect 194 1703 205 1706
rect 202 1603 205 1703
rect 234 1656 237 1726
rect 226 1653 237 1656
rect 210 1623 213 1636
rect 154 1573 165 1576
rect 162 1523 165 1573
rect 130 1393 133 1416
rect 90 1226 93 1256
rect 82 1223 93 1226
rect 114 1226 117 1326
rect 162 1236 165 1336
rect 170 1333 173 1546
rect 178 1503 181 1536
rect 218 1513 221 1616
rect 226 1603 229 1653
rect 234 1586 237 1626
rect 230 1583 237 1586
rect 186 1413 197 1416
rect 218 1403 221 1506
rect 230 1446 233 1583
rect 230 1443 237 1446
rect 234 1423 237 1443
rect 226 1403 229 1416
rect 186 1333 189 1346
rect 178 1313 181 1326
rect 194 1256 197 1376
rect 218 1333 221 1396
rect 234 1356 237 1416
rect 226 1353 237 1356
rect 226 1326 229 1353
rect 242 1336 245 1636
rect 266 1623 269 1786
rect 282 1733 285 1806
rect 290 1803 293 1926
rect 322 1836 325 1926
rect 354 1906 357 1926
rect 346 1903 357 1906
rect 346 1846 349 1903
rect 346 1843 357 1846
rect 314 1833 325 1836
rect 298 1813 301 1826
rect 274 1703 277 1716
rect 282 1703 285 1716
rect 298 1646 301 1796
rect 282 1643 301 1646
rect 266 1576 269 1616
rect 258 1573 269 1576
rect 258 1533 261 1573
rect 282 1536 285 1643
rect 314 1603 317 1833
rect 330 1756 333 1826
rect 330 1753 337 1756
rect 322 1713 325 1736
rect 334 1706 337 1753
rect 330 1703 337 1706
rect 346 1703 349 1816
rect 354 1783 357 1843
rect 362 1813 365 1946
rect 514 1943 517 1966
rect 362 1733 365 1796
rect 370 1776 373 1826
rect 378 1793 381 1806
rect 386 1783 389 1796
rect 370 1773 377 1776
rect 374 1706 377 1773
rect 394 1733 397 1926
rect 434 1923 437 1936
rect 538 1933 541 1946
rect 450 1906 453 1926
rect 442 1903 453 1906
rect 410 1813 413 1826
rect 442 1793 445 1903
rect 474 1803 477 1926
rect 538 1856 541 1916
rect 554 1896 557 1926
rect 570 1896 573 1966
rect 618 1933 621 1946
rect 554 1893 565 1896
rect 570 1893 581 1896
rect 538 1853 549 1856
rect 522 1793 525 1816
rect 546 1776 549 1853
rect 562 1823 565 1893
rect 578 1836 581 1893
rect 626 1836 629 1956
rect 730 1953 733 2040
rect 978 1956 981 1976
rect 978 1953 985 1956
rect 570 1833 581 1836
rect 610 1833 629 1836
rect 698 1926 701 1946
rect 714 1933 733 1936
rect 698 1923 709 1926
rect 570 1816 573 1833
rect 562 1813 573 1816
rect 562 1793 565 1806
rect 538 1773 549 1776
rect 370 1703 377 1706
rect 330 1623 333 1703
rect 370 1686 373 1703
rect 362 1683 373 1686
rect 362 1626 365 1683
rect 386 1636 389 1716
rect 378 1633 389 1636
rect 362 1623 373 1626
rect 370 1603 373 1623
rect 378 1613 381 1633
rect 426 1613 429 1736
rect 458 1733 461 1746
rect 474 1716 477 1736
rect 482 1733 485 1746
rect 434 1703 437 1716
rect 466 1713 477 1716
rect 466 1636 469 1713
rect 466 1633 477 1636
rect 266 1533 285 1536
rect 354 1543 381 1546
rect 394 1543 397 1606
rect 250 1373 253 1526
rect 258 1403 261 1426
rect 242 1333 253 1336
rect 266 1333 269 1533
rect 282 1506 285 1526
rect 282 1503 293 1506
rect 346 1503 349 1526
rect 290 1436 293 1503
rect 282 1433 293 1436
rect 282 1413 285 1433
rect 194 1253 205 1256
rect 154 1233 165 1236
rect 114 1223 125 1226
rect 82 1133 85 1223
rect 98 1123 101 1216
rect 122 1176 125 1223
rect 114 1173 125 1176
rect 114 1133 117 1173
rect 138 1113 141 1156
rect 146 1136 149 1216
rect 154 1203 157 1233
rect 202 1203 205 1253
rect 210 1233 213 1326
rect 218 1323 229 1326
rect 218 1313 221 1323
rect 234 1313 237 1326
rect 242 1253 245 1326
rect 250 1246 253 1333
rect 274 1323 277 1336
rect 234 1243 253 1246
rect 234 1226 237 1243
rect 210 1223 237 1226
rect 210 1153 213 1223
rect 226 1203 229 1216
rect 234 1143 237 1206
rect 250 1196 253 1236
rect 258 1205 261 1256
rect 314 1236 317 1346
rect 322 1306 325 1336
rect 338 1313 341 1406
rect 354 1403 357 1543
rect 370 1413 381 1416
rect 402 1413 405 1526
rect 434 1516 437 1546
rect 442 1543 445 1576
rect 474 1573 477 1633
rect 482 1613 485 1706
rect 498 1623 501 1636
rect 538 1613 541 1773
rect 554 1723 557 1736
rect 578 1713 581 1726
rect 482 1563 485 1606
rect 498 1593 509 1596
rect 450 1533 453 1546
rect 498 1533 501 1593
rect 434 1513 445 1516
rect 498 1513 501 1526
rect 506 1523 509 1546
rect 522 1513 525 1566
rect 426 1423 429 1436
rect 410 1403 413 1416
rect 370 1323 381 1326
rect 322 1303 349 1306
rect 370 1303 373 1316
rect 386 1306 389 1386
rect 418 1383 421 1416
rect 402 1333 413 1336
rect 426 1333 429 1366
rect 394 1313 397 1326
rect 402 1306 405 1316
rect 386 1303 405 1306
rect 410 1296 413 1333
rect 418 1303 421 1326
rect 314 1233 325 1236
rect 266 1213 269 1226
rect 282 1213 293 1216
rect 314 1213 317 1226
rect 266 1196 269 1206
rect 250 1193 269 1196
rect 146 1133 165 1136
rect 162 1036 165 1126
rect 170 1056 173 1136
rect 218 1113 221 1136
rect 234 1103 237 1136
rect 258 1123 261 1146
rect 314 1123 317 1206
rect 322 1205 325 1233
rect 338 1213 341 1296
rect 394 1293 413 1296
rect 394 1213 397 1293
rect 402 1133 405 1146
rect 170 1053 189 1056
rect 154 1033 165 1036
rect 154 1003 157 1033
rect 178 1013 181 1036
rect 186 1013 189 1053
rect 226 1013 229 1026
rect 82 613 85 806
rect 98 763 101 816
rect 122 753 125 946
rect 154 903 157 926
rect 170 913 173 936
rect 178 933 181 946
rect 186 913 189 926
rect 202 923 205 1006
rect 210 843 213 956
rect 234 953 237 1006
rect 242 993 245 1006
rect 250 996 253 1026
rect 282 1013 285 1026
rect 306 1003 309 1026
rect 322 1013 325 1026
rect 338 1013 341 1126
rect 354 1113 357 1126
rect 410 1113 413 1126
rect 418 1103 421 1216
rect 442 1213 445 1513
rect 450 1413 453 1426
rect 482 1403 485 1436
rect 490 1323 493 1346
rect 530 1333 533 1526
rect 546 1433 549 1536
rect 562 1523 565 1616
rect 546 1366 549 1416
rect 554 1413 557 1426
rect 538 1363 549 1366
rect 538 1316 541 1363
rect 546 1333 549 1346
rect 546 1323 565 1326
rect 538 1313 549 1316
rect 570 1283 573 1366
rect 578 1313 581 1606
rect 586 1603 589 1806
rect 610 1746 613 1833
rect 650 1803 653 1816
rect 610 1743 621 1746
rect 618 1643 621 1743
rect 634 1703 637 1796
rect 666 1793 669 1806
rect 642 1723 661 1726
rect 626 1623 629 1636
rect 642 1613 645 1723
rect 650 1703 653 1716
rect 650 1613 653 1636
rect 658 1613 661 1626
rect 682 1623 685 1806
rect 698 1803 701 1923
rect 706 1606 709 1746
rect 714 1723 717 1736
rect 730 1723 733 1933
rect 778 1923 781 1946
rect 802 1923 805 1936
rect 818 1933 821 1946
rect 770 1753 773 1816
rect 818 1813 821 1916
rect 842 1806 845 1936
rect 778 1793 781 1806
rect 786 1733 789 1806
rect 818 1803 845 1806
rect 874 1803 877 1936
rect 914 1846 917 1936
rect 906 1843 917 1846
rect 882 1813 885 1836
rect 818 1746 821 1803
rect 898 1796 901 1806
rect 818 1743 829 1746
rect 794 1726 797 1736
rect 602 1503 605 1536
rect 626 1523 629 1606
rect 642 1603 653 1606
rect 650 1593 653 1603
rect 690 1603 709 1606
rect 754 1603 757 1726
rect 770 1713 773 1726
rect 794 1723 805 1726
rect 794 1693 797 1716
rect 802 1613 805 1723
rect 810 1703 813 1726
rect 690 1523 693 1603
rect 698 1533 701 1596
rect 474 1143 477 1216
rect 490 1133 493 1156
rect 250 993 261 996
rect 258 933 261 993
rect 234 913 237 926
rect 186 813 189 836
rect 154 793 157 806
rect 202 803 205 826
rect 218 813 221 826
rect 226 806 229 836
rect 234 813 237 846
rect 210 793 213 806
rect 226 803 237 806
rect 130 653 133 766
rect 146 713 149 726
rect 154 723 157 756
rect 170 723 173 746
rect 178 716 181 736
rect 234 733 237 803
rect 258 723 261 806
rect 266 743 269 936
rect 290 813 293 826
rect 298 813 301 926
rect 314 923 317 1006
rect 354 976 357 1006
rect 346 973 357 976
rect 322 913 325 936
rect 346 926 349 973
rect 362 933 365 946
rect 378 933 381 1016
rect 434 943 437 1016
rect 346 923 357 926
rect 378 923 397 926
rect 322 803 325 816
rect 354 766 357 923
rect 378 913 397 916
rect 346 763 357 766
rect 82 323 85 596
rect 106 503 109 616
rect 154 613 157 626
rect 170 616 173 716
rect 178 713 185 716
rect 182 646 185 713
rect 178 643 185 646
rect 178 623 181 643
rect 170 613 189 616
rect 210 613 213 626
rect 250 613 269 616
rect 274 613 277 736
rect 282 713 285 726
rect 298 723 301 746
rect 298 613 301 656
rect 306 613 309 726
rect 114 593 117 606
rect 178 556 181 606
rect 234 593 237 606
rect 242 603 261 606
rect 162 553 181 556
rect 162 506 165 553
rect 170 513 173 536
rect 130 403 133 506
rect 162 503 181 506
rect 194 503 197 526
rect 226 503 229 536
rect 146 413 165 416
rect 178 413 181 503
rect 234 426 237 536
rect 242 493 245 526
rect 258 513 261 603
rect 266 503 269 613
rect 330 593 333 606
rect 322 523 325 546
rect 234 423 245 426
rect 74 203 77 236
rect 114 233 117 326
rect 122 316 125 336
rect 122 313 129 316
rect 126 246 129 313
rect 138 263 141 406
rect 186 393 189 406
rect 234 403 237 416
rect 146 333 149 346
rect 170 313 173 326
rect 202 323 205 346
rect 210 333 213 366
rect 242 343 245 423
rect 258 413 261 436
rect 266 363 269 496
rect 322 413 325 426
rect 122 243 129 246
rect 98 213 101 226
rect 122 153 125 243
rect 130 146 133 226
rect 154 213 157 306
rect 122 133 125 146
rect 130 143 141 146
rect 138 123 141 143
rect 154 123 157 186
rect 162 123 165 156
rect 178 143 181 206
rect 186 183 189 266
rect 202 196 205 216
rect 210 203 213 226
rect 234 223 237 326
rect 250 303 253 326
rect 258 203 261 336
rect 202 193 213 196
rect 202 133 205 156
rect 210 126 213 193
rect 266 173 269 226
rect 322 193 325 216
rect 346 203 349 763
rect 370 753 373 806
rect 386 803 389 856
rect 394 813 397 913
rect 418 903 421 926
rect 362 723 365 746
rect 386 733 389 796
rect 410 756 413 836
rect 410 753 417 756
rect 402 733 405 746
rect 402 676 405 716
rect 394 673 405 676
rect 370 586 373 616
rect 378 613 381 626
rect 394 613 397 673
rect 414 636 417 753
rect 410 633 417 636
rect 402 606 405 626
rect 410 613 413 633
rect 426 623 429 936
rect 434 713 437 806
rect 442 803 445 1116
rect 458 933 461 1016
rect 466 1006 469 1126
rect 482 1013 485 1036
rect 466 1003 485 1006
rect 490 996 493 1026
rect 506 1013 509 1136
rect 530 1133 533 1216
rect 546 1133 549 1146
rect 514 1123 533 1126
rect 538 1123 549 1126
rect 530 1013 533 1116
rect 538 1006 541 1026
rect 442 723 445 736
rect 370 583 381 586
rect 386 583 389 606
rect 394 603 405 606
rect 362 533 365 546
rect 378 523 381 583
rect 362 503 365 516
rect 386 433 389 526
rect 362 403 365 426
rect 370 393 373 426
rect 378 303 381 416
rect 394 406 397 603
rect 402 413 405 586
rect 410 503 413 526
rect 426 496 429 616
rect 442 533 445 616
rect 450 583 453 856
rect 466 853 469 996
rect 474 993 493 996
rect 498 993 501 1006
rect 530 1003 541 1006
rect 530 996 533 1003
rect 522 993 533 996
rect 474 923 477 993
rect 482 916 485 936
rect 474 913 485 916
rect 474 813 477 913
rect 490 833 493 986
rect 522 923 525 993
rect 546 983 549 1016
rect 562 1013 565 1206
rect 586 1193 589 1326
rect 626 1323 629 1406
rect 658 1323 661 1436
rect 698 1413 701 1526
rect 706 1386 709 1406
rect 730 1393 733 1506
rect 754 1413 757 1536
rect 770 1503 773 1606
rect 802 1426 805 1596
rect 818 1593 821 1743
rect 798 1423 805 1426
rect 698 1383 709 1386
rect 690 1333 693 1346
rect 698 1343 701 1383
rect 798 1376 801 1423
rect 810 1383 813 1416
rect 826 1413 829 1516
rect 834 1513 837 1646
rect 842 1516 845 1796
rect 890 1793 901 1796
rect 906 1793 909 1843
rect 914 1823 917 1836
rect 922 1813 925 1866
rect 938 1816 941 1926
rect 954 1816 957 1946
rect 982 1886 985 1953
rect 1002 1943 1005 2040
rect 1034 2026 1037 2040
rect 1026 2023 1037 2026
rect 1026 1956 1029 2023
rect 1026 1953 1037 1956
rect 1050 1953 1053 2040
rect 1066 1973 1069 2040
rect 1138 2026 1141 2040
rect 1130 2023 1141 2026
rect 1130 1976 1133 2023
rect 1130 1973 1141 1976
rect 994 1933 1013 1936
rect 994 1923 997 1933
rect 978 1883 985 1886
rect 930 1813 941 1816
rect 946 1813 957 1816
rect 962 1813 965 1826
rect 978 1813 981 1883
rect 1002 1823 1005 1926
rect 1018 1863 1021 1926
rect 1034 1856 1037 1953
rect 1042 1923 1045 1936
rect 1026 1853 1037 1856
rect 1026 1836 1029 1853
rect 1022 1833 1029 1836
rect 930 1803 933 1813
rect 898 1746 901 1793
rect 938 1786 941 1806
rect 934 1783 941 1786
rect 898 1743 925 1746
rect 850 1716 853 1736
rect 850 1713 861 1716
rect 858 1646 861 1713
rect 898 1693 901 1726
rect 850 1643 861 1646
rect 850 1593 853 1643
rect 858 1613 861 1626
rect 906 1613 909 1736
rect 922 1713 925 1743
rect 934 1646 937 1783
rect 934 1643 941 1646
rect 874 1526 877 1606
rect 890 1593 893 1606
rect 874 1523 917 1526
rect 842 1513 853 1516
rect 850 1466 853 1513
rect 842 1463 853 1466
rect 834 1413 837 1426
rect 818 1403 837 1406
rect 798 1373 805 1376
rect 802 1353 805 1373
rect 610 1203 613 1316
rect 618 1303 621 1316
rect 626 1216 629 1266
rect 626 1213 637 1216
rect 642 1213 645 1316
rect 706 1303 709 1326
rect 674 1193 677 1286
rect 730 1223 733 1236
rect 578 1116 581 1136
rect 658 1133 661 1156
rect 578 1113 589 1116
rect 586 1026 589 1113
rect 578 1023 589 1026
rect 626 1023 629 1126
rect 674 1113 677 1136
rect 706 1123 709 1206
rect 738 1126 741 1336
rect 754 1313 757 1336
rect 778 1333 781 1346
rect 826 1333 829 1386
rect 754 1213 757 1226
rect 786 1213 789 1236
rect 794 1203 797 1316
rect 802 1306 805 1326
rect 834 1323 837 1403
rect 842 1366 845 1463
rect 858 1393 861 1406
rect 842 1363 861 1366
rect 802 1303 809 1306
rect 806 1216 809 1303
rect 834 1263 837 1316
rect 858 1256 861 1363
rect 882 1336 885 1416
rect 842 1253 861 1256
rect 874 1333 885 1336
rect 802 1213 809 1216
rect 818 1213 821 1226
rect 794 1166 797 1196
rect 786 1163 797 1166
rect 786 1143 789 1163
rect 802 1143 805 1213
rect 738 1123 757 1126
rect 554 953 557 996
rect 530 906 533 936
rect 530 903 541 906
rect 538 813 541 903
rect 578 813 581 1023
rect 602 933 605 1006
rect 626 1003 629 1016
rect 746 993 749 1116
rect 762 1103 765 1126
rect 458 783 461 806
rect 506 776 509 806
rect 602 803 605 816
rect 618 806 621 926
rect 666 833 669 926
rect 674 923 685 926
rect 690 883 693 926
rect 730 893 733 936
rect 610 803 621 806
rect 514 783 517 796
rect 498 773 509 776
rect 474 743 477 756
rect 466 603 469 646
rect 482 613 485 746
rect 498 723 501 773
rect 546 763 549 796
rect 506 733 509 746
rect 554 733 557 756
rect 506 593 509 726
rect 538 713 541 726
rect 530 603 533 626
rect 562 613 565 736
rect 610 643 613 726
rect 626 723 629 796
rect 594 613 605 616
rect 546 603 573 606
rect 530 583 533 596
rect 458 523 461 556
rect 394 403 405 406
rect 394 323 397 396
rect 402 316 405 403
rect 410 363 413 496
rect 426 493 437 496
rect 410 333 413 356
rect 434 346 437 493
rect 482 403 485 526
rect 426 343 437 346
rect 386 313 405 316
rect 362 223 365 236
rect 362 193 365 206
rect 194 123 213 126
rect 250 113 253 126
rect 274 103 277 156
rect 282 123 285 146
rect 330 133 333 146
rect 338 133 341 176
rect 298 113 301 126
rect 346 123 349 156
rect 378 153 381 216
rect 386 213 389 313
rect 394 156 397 216
rect 402 193 405 306
rect 410 213 413 236
rect 426 213 429 343
rect 442 313 445 326
rect 490 323 493 426
rect 538 416 541 526
rect 546 523 549 603
rect 618 593 621 606
rect 634 603 637 806
rect 642 733 645 826
rect 738 823 741 936
rect 770 933 773 1136
rect 786 1133 805 1136
rect 786 1123 789 1133
rect 802 1113 805 1126
rect 810 1123 813 1196
rect 842 1183 845 1253
rect 874 1236 877 1333
rect 874 1233 885 1236
rect 882 1213 885 1233
rect 842 1133 845 1146
rect 858 1123 861 1206
rect 874 1133 877 1146
rect 778 933 781 1106
rect 786 933 789 1016
rect 754 913 757 926
rect 770 923 781 926
rect 810 923 813 946
rect 786 833 789 916
rect 650 813 669 816
rect 682 813 693 816
rect 770 813 789 816
rect 650 803 653 813
rect 794 803 797 896
rect 826 803 829 856
rect 834 803 837 936
rect 866 933 869 1016
rect 874 1013 877 1026
rect 882 1003 885 1146
rect 890 1123 893 1326
rect 898 1303 901 1506
rect 906 1393 909 1416
rect 914 1326 917 1336
rect 906 1323 917 1326
rect 906 1286 909 1323
rect 902 1283 909 1286
rect 902 1196 905 1283
rect 914 1203 917 1316
rect 922 1306 925 1586
rect 930 1406 933 1516
rect 938 1413 941 1643
rect 946 1613 949 1813
rect 946 1523 949 1606
rect 954 1583 957 1806
rect 978 1793 981 1806
rect 962 1623 965 1736
rect 1010 1733 1013 1816
rect 1022 1776 1025 1833
rect 1050 1813 1069 1816
rect 1090 1813 1093 1936
rect 1098 1923 1101 1946
rect 1106 1906 1109 1936
rect 1102 1903 1109 1906
rect 1102 1826 1105 1903
rect 1098 1823 1105 1826
rect 1022 1773 1029 1776
rect 930 1403 949 1406
rect 946 1323 949 1346
rect 954 1333 957 1416
rect 962 1386 965 1536
rect 986 1533 989 1546
rect 986 1496 989 1516
rect 978 1493 989 1496
rect 978 1436 981 1493
rect 978 1433 989 1436
rect 986 1413 989 1433
rect 970 1393 973 1406
rect 994 1403 997 1616
rect 1002 1613 1005 1716
rect 1018 1603 1021 1656
rect 1026 1633 1029 1773
rect 1042 1733 1045 1746
rect 1050 1653 1053 1813
rect 1066 1793 1069 1813
rect 1074 1603 1077 1806
rect 1026 1523 1029 1546
rect 1010 1413 1013 1426
rect 1026 1423 1029 1436
rect 1034 1423 1037 1446
rect 1026 1403 1029 1416
rect 962 1383 981 1386
rect 962 1343 965 1383
rect 1042 1343 1045 1586
rect 1074 1533 1077 1546
rect 1050 1413 1053 1436
rect 1058 1333 1061 1406
rect 954 1313 957 1326
rect 922 1303 933 1306
rect 930 1236 933 1303
rect 1018 1296 1021 1316
rect 1026 1296 1029 1306
rect 1018 1293 1029 1296
rect 922 1233 933 1236
rect 902 1193 909 1196
rect 922 1193 925 1233
rect 946 1213 965 1216
rect 1018 1206 1021 1226
rect 1026 1223 1029 1293
rect 906 1176 909 1193
rect 906 1173 917 1176
rect 914 1116 917 1173
rect 906 1113 917 1116
rect 906 1023 909 1113
rect 922 1013 925 1026
rect 906 993 909 1006
rect 938 1005 941 1016
rect 962 1013 965 1206
rect 1018 1203 1037 1206
rect 1050 1203 1053 1326
rect 1066 1313 1069 1416
rect 1066 1213 1069 1306
rect 1034 1133 1037 1203
rect 1058 1133 1061 1206
rect 1026 1116 1029 1126
rect 1034 1116 1037 1126
rect 1074 1123 1077 1436
rect 1082 1366 1085 1446
rect 1090 1383 1093 1406
rect 1082 1363 1089 1366
rect 1086 1286 1089 1363
rect 1082 1283 1089 1286
rect 1098 1283 1101 1823
rect 1114 1323 1117 1956
rect 1138 1933 1141 1973
rect 1154 1953 1157 2040
rect 1130 1806 1133 1926
rect 1138 1913 1141 1926
rect 1154 1866 1157 1926
rect 1154 1863 1165 1866
rect 1126 1803 1133 1806
rect 1126 1746 1129 1803
rect 1126 1743 1133 1746
rect 1122 1713 1125 1726
rect 1130 1723 1133 1743
rect 1138 1543 1141 1796
rect 1146 1733 1149 1826
rect 1154 1783 1157 1836
rect 1162 1786 1165 1863
rect 1170 1803 1173 1926
rect 1178 1813 1181 1826
rect 1186 1806 1189 1936
rect 1202 1933 1213 1936
rect 1202 1833 1205 1933
rect 1178 1803 1189 1806
rect 1162 1783 1169 1786
rect 1154 1703 1157 1736
rect 1166 1696 1169 1783
rect 1178 1743 1181 1803
rect 1194 1713 1197 1816
rect 1210 1783 1213 1806
rect 1218 1726 1221 1966
rect 1258 1963 1261 2040
rect 1234 1933 1237 1946
rect 1234 1823 1237 1916
rect 1250 1866 1253 1936
rect 1274 1923 1277 1946
rect 1242 1863 1253 1866
rect 1226 1793 1229 1806
rect 1234 1733 1237 1806
rect 1242 1793 1245 1863
rect 1242 1733 1245 1746
rect 1202 1713 1205 1726
rect 1218 1723 1229 1726
rect 1162 1693 1169 1696
rect 1162 1646 1165 1693
rect 1226 1646 1229 1723
rect 1162 1643 1173 1646
rect 1226 1643 1237 1646
rect 1170 1576 1173 1643
rect 1146 1573 1173 1576
rect 1130 1416 1133 1536
rect 1126 1413 1133 1416
rect 1126 1366 1129 1413
rect 1126 1363 1133 1366
rect 1130 1346 1133 1363
rect 1138 1353 1141 1406
rect 1130 1343 1141 1346
rect 1130 1323 1133 1336
rect 1138 1293 1141 1343
rect 1146 1323 1149 1573
rect 1186 1533 1189 1616
rect 1218 1546 1221 1616
rect 1226 1613 1229 1626
rect 1210 1543 1221 1546
rect 1154 1506 1157 1526
rect 1210 1516 1213 1543
rect 1202 1513 1213 1516
rect 1154 1503 1165 1506
rect 1162 1446 1165 1503
rect 1154 1443 1165 1446
rect 1202 1446 1205 1513
rect 1202 1443 1213 1446
rect 1154 1303 1157 1443
rect 1162 1333 1165 1426
rect 1178 1323 1181 1406
rect 1210 1363 1213 1443
rect 1218 1403 1221 1516
rect 1234 1406 1237 1643
rect 1250 1613 1253 1856
rect 1282 1853 1285 2040
rect 1298 2026 1301 2040
rect 1298 2023 1309 2026
rect 1306 1976 1309 2023
rect 1298 1973 1309 1976
rect 1298 1956 1301 1973
rect 1294 1953 1301 1956
rect 1294 1886 1297 1953
rect 1330 1943 1341 1946
rect 1330 1893 1333 1943
rect 1346 1936 1349 2040
rect 1434 1946 1437 2040
rect 1482 1946 1485 2040
rect 1338 1913 1341 1936
rect 1346 1933 1357 1936
rect 1378 1933 1381 1946
rect 1426 1943 1437 1946
rect 1466 1943 1485 1946
rect 1490 1943 1509 1946
rect 1294 1883 1301 1886
rect 1258 1766 1261 1816
rect 1258 1763 1269 1766
rect 1266 1646 1269 1763
rect 1282 1723 1285 1736
rect 1258 1643 1269 1646
rect 1250 1593 1253 1606
rect 1258 1603 1261 1643
rect 1290 1633 1293 1736
rect 1298 1716 1301 1883
rect 1314 1733 1317 1816
rect 1338 1793 1341 1806
rect 1354 1786 1357 1933
rect 1370 1813 1373 1826
rect 1346 1783 1357 1786
rect 1298 1713 1309 1716
rect 1306 1636 1309 1713
rect 1306 1633 1325 1636
rect 1242 1513 1245 1526
rect 1266 1523 1269 1616
rect 1282 1613 1285 1626
rect 1314 1546 1317 1606
rect 1322 1573 1325 1633
rect 1306 1543 1317 1546
rect 1306 1523 1309 1543
rect 1250 1413 1253 1436
rect 1234 1403 1245 1406
rect 1242 1346 1245 1403
rect 1226 1333 1229 1346
rect 1242 1343 1261 1346
rect 1250 1323 1253 1336
rect 1258 1333 1261 1343
rect 1258 1293 1261 1326
rect 1266 1323 1269 1406
rect 1274 1323 1277 1516
rect 1314 1513 1317 1526
rect 1298 1493 1301 1506
rect 1322 1503 1325 1526
rect 1282 1303 1285 1426
rect 1346 1403 1349 1783
rect 1394 1776 1397 1826
rect 1410 1803 1413 1926
rect 1426 1896 1429 1943
rect 1434 1923 1437 1936
rect 1422 1893 1429 1896
rect 1422 1816 1425 1893
rect 1422 1813 1429 1816
rect 1434 1813 1437 1916
rect 1394 1773 1405 1776
rect 1386 1696 1389 1716
rect 1378 1693 1389 1696
rect 1378 1646 1381 1693
rect 1378 1643 1389 1646
rect 1378 1603 1381 1626
rect 1386 1613 1389 1643
rect 1394 1606 1397 1766
rect 1402 1646 1405 1773
rect 1402 1643 1413 1646
rect 1402 1623 1405 1643
rect 1386 1603 1397 1606
rect 1362 1493 1365 1526
rect 1370 1476 1373 1536
rect 1362 1473 1373 1476
rect 1362 1366 1365 1473
rect 1290 1333 1293 1366
rect 1362 1363 1373 1366
rect 1082 1203 1085 1283
rect 1146 1206 1149 1286
rect 1314 1226 1317 1246
rect 1178 1223 1197 1226
rect 1178 1213 1181 1223
rect 1186 1206 1189 1216
rect 1194 1213 1197 1223
rect 1306 1223 1317 1226
rect 1106 1123 1109 1206
rect 1138 1193 1141 1206
rect 1146 1203 1173 1206
rect 1186 1203 1197 1206
rect 1170 1173 1173 1203
rect 1170 1133 1173 1166
rect 1178 1133 1181 1196
rect 1194 1193 1197 1203
rect 1226 1133 1229 1176
rect 1018 1113 1037 1116
rect 1018 1013 1021 1113
rect 1018 966 1021 996
rect 1034 993 1037 1006
rect 1010 963 1021 966
rect 954 916 957 936
rect 850 813 853 836
rect 866 813 869 916
rect 946 913 957 916
rect 946 826 949 913
rect 946 823 957 826
rect 850 803 861 806
rect 954 803 957 823
rect 962 803 965 816
rect 970 813 973 926
rect 978 906 981 936
rect 978 903 989 906
rect 986 836 989 903
rect 978 833 989 836
rect 1010 836 1013 963
rect 1026 933 1029 946
rect 1058 933 1061 1016
rect 1114 1003 1117 1016
rect 1122 1013 1125 1026
rect 1130 986 1133 1126
rect 1234 1103 1237 1126
rect 1114 983 1133 986
rect 1010 833 1021 836
rect 978 803 981 833
rect 994 793 997 806
rect 658 746 661 766
rect 650 646 653 746
rect 658 743 677 746
rect 646 643 653 646
rect 646 566 649 643
rect 674 636 677 743
rect 778 733 789 736
rect 746 713 749 726
rect 658 633 677 636
rect 646 563 653 566
rect 562 543 573 546
rect 562 493 565 543
rect 530 413 541 416
rect 578 413 581 536
rect 626 533 629 546
rect 650 543 653 563
rect 602 496 605 526
rect 594 493 605 496
rect 594 416 597 493
rect 594 413 605 416
rect 506 403 517 406
rect 530 326 533 413
rect 514 323 533 326
rect 394 153 413 156
rect 402 133 405 146
rect 354 113 357 126
rect 378 113 381 126
rect 402 103 405 126
rect 410 113 413 153
rect 466 133 469 146
rect 474 126 477 216
rect 498 203 501 246
rect 514 236 517 323
rect 538 243 541 326
rect 506 233 517 236
rect 506 203 509 233
rect 554 203 557 336
rect 562 296 565 366
rect 602 363 605 413
rect 610 353 613 526
rect 626 506 629 526
rect 658 523 661 633
rect 626 503 637 506
rect 634 446 637 503
rect 626 443 637 446
rect 618 333 621 406
rect 626 346 629 443
rect 674 436 677 616
rect 682 613 693 616
rect 690 523 693 546
rect 698 513 701 656
rect 738 616 741 636
rect 754 616 757 726
rect 770 703 773 726
rect 786 633 789 726
rect 802 693 805 726
rect 810 623 813 736
rect 850 733 853 746
rect 842 623 845 726
rect 858 713 861 726
rect 730 613 741 616
rect 750 613 757 616
rect 730 556 733 613
rect 750 566 753 613
rect 746 563 753 566
rect 730 553 741 556
rect 674 433 693 436
rect 634 393 637 406
rect 626 343 653 346
rect 674 343 677 386
rect 634 296 637 326
rect 562 293 573 296
rect 570 226 573 293
rect 626 293 637 296
rect 626 236 629 293
rect 650 266 653 343
rect 682 333 685 406
rect 690 376 693 433
rect 706 393 709 546
rect 714 523 717 536
rect 730 506 733 526
rect 722 503 733 506
rect 722 426 725 503
rect 722 423 733 426
rect 730 403 733 423
rect 738 396 741 553
rect 746 476 749 563
rect 762 513 765 606
rect 858 583 861 616
rect 874 613 877 726
rect 962 723 965 746
rect 970 743 973 756
rect 890 613 893 626
rect 810 533 813 556
rect 746 473 757 476
rect 730 393 741 396
rect 730 376 733 393
rect 690 373 701 376
rect 698 326 701 373
rect 642 263 653 266
rect 690 323 701 326
rect 722 373 733 376
rect 626 233 637 236
rect 562 223 573 226
rect 562 173 565 223
rect 570 193 573 206
rect 530 133 533 146
rect 458 123 477 126
rect 506 113 509 126
rect 538 123 541 136
rect 570 133 573 156
rect 554 113 557 126
rect 578 113 581 136
rect 586 123 589 216
rect 634 213 637 233
rect 642 203 645 263
rect 650 213 653 226
rect 658 213 661 246
rect 642 133 645 156
rect 674 123 677 146
rect 690 116 693 323
rect 722 236 725 373
rect 754 366 757 473
rect 786 413 789 526
rect 826 513 829 526
rect 882 523 885 606
rect 962 603 965 636
rect 970 603 973 736
rect 986 706 989 736
rect 1002 723 1005 816
rect 1018 796 1021 833
rect 1034 813 1037 926
rect 1058 913 1061 926
rect 1066 903 1069 916
rect 1114 856 1117 983
rect 1138 863 1141 1016
rect 1146 1013 1149 1026
rect 1178 1013 1181 1056
rect 1242 1053 1245 1136
rect 1282 1033 1285 1196
rect 1306 1166 1309 1223
rect 1306 1163 1317 1166
rect 1314 1143 1317 1163
rect 1322 1156 1325 1206
rect 1330 1163 1333 1326
rect 1338 1243 1341 1326
rect 1362 1323 1365 1336
rect 1370 1333 1373 1363
rect 1378 1303 1381 1536
rect 1386 1516 1389 1603
rect 1410 1536 1413 1626
rect 1418 1613 1421 1796
rect 1426 1763 1429 1813
rect 1450 1723 1453 1936
rect 1466 1876 1469 1943
rect 1482 1883 1485 1936
rect 1490 1886 1493 1943
rect 1514 1933 1517 1946
rect 1498 1903 1501 1926
rect 1554 1923 1557 1946
rect 1658 1933 1661 1946
rect 1666 1943 1669 1956
rect 1722 1936 1725 1956
rect 1722 1933 1733 1936
rect 1810 1933 1813 1946
rect 1578 1923 1589 1926
rect 1490 1883 1501 1886
rect 1466 1873 1477 1876
rect 1474 1766 1477 1873
rect 1466 1763 1477 1766
rect 1466 1726 1469 1763
rect 1458 1723 1469 1726
rect 1498 1723 1501 1883
rect 1546 1803 1549 1916
rect 1570 1803 1573 1906
rect 1578 1903 1581 1916
rect 1642 1803 1645 1926
rect 1562 1783 1565 1796
rect 1394 1533 1413 1536
rect 1450 1516 1453 1536
rect 1458 1523 1461 1723
rect 1514 1676 1517 1736
rect 1514 1673 1533 1676
rect 1466 1623 1493 1626
rect 1466 1613 1469 1623
rect 1466 1533 1469 1606
rect 1474 1593 1477 1616
rect 1386 1513 1397 1516
rect 1394 1446 1397 1513
rect 1386 1443 1397 1446
rect 1442 1513 1453 1516
rect 1386 1326 1389 1443
rect 1442 1436 1445 1513
rect 1442 1433 1453 1436
rect 1466 1433 1469 1526
rect 1394 1333 1397 1426
rect 1410 1413 1429 1416
rect 1410 1403 1437 1406
rect 1410 1333 1413 1346
rect 1386 1323 1397 1326
rect 1434 1323 1437 1403
rect 1450 1353 1453 1433
rect 1474 1413 1477 1426
rect 1466 1363 1469 1406
rect 1482 1346 1485 1526
rect 1490 1423 1493 1606
rect 1506 1533 1509 1616
rect 1530 1583 1533 1673
rect 1538 1593 1541 1616
rect 1554 1613 1557 1726
rect 1586 1613 1589 1796
rect 1610 1736 1613 1786
rect 1650 1753 1653 1806
rect 1594 1733 1613 1736
rect 1666 1733 1669 1816
rect 1674 1813 1677 1926
rect 1682 1803 1685 1816
rect 1714 1803 1717 1886
rect 1722 1873 1725 1926
rect 1730 1813 1733 1933
rect 1762 1886 1765 1926
rect 1754 1883 1765 1886
rect 1826 1883 1829 1936
rect 1674 1733 1677 1756
rect 1594 1723 1597 1733
rect 1594 1613 1597 1636
rect 1602 1613 1605 1726
rect 1634 1623 1637 1646
rect 1594 1596 1597 1606
rect 1618 1603 1621 1616
rect 1650 1603 1653 1726
rect 1722 1696 1725 1736
rect 1714 1693 1725 1696
rect 1730 1696 1733 1806
rect 1754 1803 1757 1883
rect 1762 1803 1765 1876
rect 1770 1706 1773 1726
rect 1762 1703 1773 1706
rect 1730 1693 1741 1696
rect 1714 1603 1717 1693
rect 1594 1593 1605 1596
rect 1498 1496 1501 1526
rect 1506 1513 1509 1526
rect 1498 1493 1509 1496
rect 1506 1436 1509 1493
rect 1594 1436 1597 1586
rect 1602 1576 1605 1593
rect 1602 1573 1621 1576
rect 1498 1433 1509 1436
rect 1578 1433 1597 1436
rect 1498 1413 1501 1433
rect 1530 1413 1533 1426
rect 1474 1343 1485 1346
rect 1338 1173 1341 1216
rect 1322 1153 1341 1156
rect 1298 1133 1333 1136
rect 1290 1113 1293 1126
rect 1306 1103 1309 1126
rect 1314 1043 1317 1126
rect 1306 1013 1309 1026
rect 1194 993 1197 1006
rect 1202 976 1205 1006
rect 1198 973 1205 976
rect 1170 923 1173 936
rect 1178 903 1181 926
rect 1114 853 1133 856
rect 1186 853 1189 936
rect 1090 813 1093 826
rect 1018 793 1029 796
rect 1090 793 1093 806
rect 1026 716 1029 793
rect 1090 733 1093 746
rect 1098 733 1101 756
rect 1018 713 1029 716
rect 986 703 997 706
rect 994 636 997 703
rect 986 633 997 636
rect 986 613 989 633
rect 1018 553 1021 713
rect 1114 653 1117 816
rect 1130 803 1133 853
rect 1198 846 1201 973
rect 1210 933 1213 1006
rect 1330 996 1333 1036
rect 1338 1003 1341 1153
rect 1346 1013 1349 1166
rect 1354 1133 1357 1216
rect 1362 1163 1365 1216
rect 1370 1213 1381 1216
rect 1394 1213 1397 1323
rect 1474 1286 1477 1343
rect 1490 1313 1493 1326
rect 1498 1323 1501 1366
rect 1506 1313 1509 1336
rect 1538 1333 1541 1356
rect 1578 1343 1581 1433
rect 1618 1366 1621 1573
rect 1650 1393 1653 1526
rect 1690 1466 1693 1556
rect 1738 1553 1741 1693
rect 1762 1646 1765 1703
rect 1762 1643 1773 1646
rect 1778 1643 1781 1826
rect 1850 1746 1853 1946
rect 1858 1933 1869 1936
rect 1882 1933 1893 1936
rect 1866 1923 1885 1926
rect 1882 1883 1885 1916
rect 1890 1876 1893 1933
rect 1882 1873 1893 1876
rect 1882 1813 1885 1873
rect 1914 1816 1917 1936
rect 1930 1933 1933 1946
rect 1978 1923 1981 1946
rect 2026 1933 2037 1936
rect 2058 1933 2061 1946
rect 1914 1813 1933 1816
rect 1938 1813 1941 1886
rect 1946 1813 1949 1826
rect 1834 1743 1853 1746
rect 1770 1623 1773 1643
rect 1794 1626 1797 1716
rect 1834 1666 1837 1743
rect 1850 1716 1853 1736
rect 1890 1733 1901 1736
rect 1850 1713 1861 1716
rect 1858 1666 1861 1713
rect 1834 1663 1845 1666
rect 1786 1623 1797 1626
rect 1770 1593 1773 1606
rect 1730 1533 1733 1546
rect 1746 1533 1749 1546
rect 1674 1463 1693 1466
rect 1602 1363 1621 1366
rect 1602 1346 1605 1363
rect 1674 1353 1677 1463
rect 1682 1413 1693 1416
rect 1698 1403 1701 1526
rect 1706 1396 1709 1426
rect 1714 1413 1717 1426
rect 1594 1343 1605 1346
rect 1546 1323 1557 1326
rect 1466 1283 1477 1286
rect 1450 1193 1453 1206
rect 1354 1106 1357 1126
rect 1354 1103 1365 1106
rect 1402 1103 1405 1136
rect 1466 1133 1469 1283
rect 1498 1236 1501 1306
rect 1490 1233 1501 1236
rect 1490 1186 1493 1233
rect 1562 1213 1565 1336
rect 1594 1326 1597 1343
rect 1586 1323 1597 1326
rect 1570 1303 1573 1316
rect 1586 1266 1589 1323
rect 1586 1263 1593 1266
rect 1590 1206 1593 1263
rect 1602 1213 1605 1336
rect 1610 1306 1613 1336
rect 1610 1303 1621 1306
rect 1618 1226 1621 1303
rect 1610 1223 1621 1226
rect 1522 1193 1525 1206
rect 1590 1203 1597 1206
rect 1610 1203 1613 1223
rect 1490 1183 1501 1186
rect 1498 1136 1501 1183
rect 1594 1143 1597 1203
rect 1650 1193 1653 1206
rect 1682 1203 1685 1396
rect 1698 1393 1709 1396
rect 1698 1323 1701 1393
rect 1706 1213 1709 1336
rect 1722 1303 1725 1316
rect 1730 1226 1733 1526
rect 1786 1523 1789 1623
rect 1802 1503 1805 1646
rect 1818 1543 1821 1606
rect 1842 1593 1845 1663
rect 1850 1663 1861 1666
rect 1850 1613 1853 1663
rect 1898 1606 1901 1616
rect 1906 1613 1909 1726
rect 1930 1713 1933 1813
rect 1970 1743 1973 1756
rect 1962 1636 1965 1736
rect 1970 1713 1973 1736
rect 1978 1723 1981 1806
rect 1986 1753 1989 1886
rect 2010 1883 2013 1926
rect 2034 1813 2037 1826
rect 2042 1813 2045 1826
rect 2042 1756 2045 1806
rect 2058 1803 2061 1826
rect 2066 1813 2069 1916
rect 2042 1753 2061 1756
rect 2034 1713 2037 1746
rect 2042 1723 2045 1736
rect 2058 1723 2061 1753
rect 1954 1633 1965 1636
rect 1898 1603 1909 1606
rect 1906 1576 1909 1603
rect 1898 1573 1909 1576
rect 1898 1543 1901 1573
rect 1810 1513 1813 1526
rect 1818 1436 1821 1526
rect 1850 1513 1853 1526
rect 1882 1496 1885 1536
rect 1874 1493 1885 1496
rect 1874 1436 1877 1493
rect 1898 1483 1901 1536
rect 1930 1526 1933 1596
rect 1954 1586 1957 1633
rect 1978 1593 1981 1606
rect 1954 1583 1973 1586
rect 1922 1523 1933 1526
rect 1802 1423 1805 1436
rect 1810 1423 1813 1436
rect 1818 1433 1829 1436
rect 1810 1413 1821 1416
rect 1826 1406 1829 1433
rect 1778 1343 1789 1346
rect 1778 1333 1781 1343
rect 1730 1223 1737 1226
rect 1722 1186 1725 1216
rect 1714 1183 1725 1186
rect 1498 1133 1509 1136
rect 1354 1013 1357 1046
rect 1362 1013 1365 1103
rect 1346 996 1349 1006
rect 1458 1003 1461 1026
rect 1466 1003 1469 1126
rect 1490 1113 1493 1126
rect 1498 1013 1501 1056
rect 1506 1033 1509 1133
rect 1570 1123 1589 1126
rect 1682 1076 1685 1126
rect 1682 1073 1689 1076
rect 1218 976 1221 996
rect 1330 993 1349 996
rect 1218 973 1229 976
rect 1198 843 1205 846
rect 1154 803 1157 826
rect 1194 813 1197 826
rect 1202 803 1205 843
rect 1210 813 1213 886
rect 1226 836 1229 973
rect 1218 833 1229 836
rect 1218 743 1221 833
rect 1050 616 1053 626
rect 1050 613 1061 616
rect 914 516 917 536
rect 954 533 965 536
rect 906 513 917 516
rect 906 446 909 513
rect 906 443 917 446
rect 746 363 757 366
rect 722 233 733 236
rect 730 216 733 233
rect 722 183 725 216
rect 730 213 737 216
rect 674 113 693 116
rect 674 0 677 113
rect 698 103 701 126
rect 722 113 725 176
rect 734 156 737 213
rect 746 173 749 363
rect 778 343 781 406
rect 842 403 853 406
rect 874 403 877 416
rect 762 163 765 206
rect 810 183 813 346
rect 818 333 821 346
rect 874 333 877 346
rect 842 243 845 326
rect 730 153 737 156
rect 730 93 733 153
rect 738 123 741 136
rect 754 0 757 116
rect 786 103 789 146
rect 794 113 797 126
rect 802 123 805 156
rect 818 143 821 216
rect 842 193 845 206
rect 826 133 829 156
rect 818 113 821 126
rect 834 113 837 136
rect 882 133 885 156
rect 858 113 861 126
rect 890 113 893 216
rect 898 203 901 266
rect 906 213 909 426
rect 914 403 917 443
rect 930 413 933 526
rect 946 383 949 516
rect 962 403 965 526
rect 994 523 997 536
rect 914 203 917 246
rect 922 213 925 226
rect 978 213 981 406
rect 1018 366 1021 416
rect 1042 413 1045 556
rect 1058 523 1061 613
rect 1130 603 1133 626
rect 1138 603 1141 716
rect 1154 526 1157 606
rect 1178 563 1181 726
rect 1218 696 1221 736
rect 1226 726 1229 816
rect 1250 793 1253 936
rect 1258 933 1261 946
rect 1314 933 1317 946
rect 1258 913 1261 926
rect 1282 913 1285 926
rect 1258 813 1261 826
rect 1290 813 1293 926
rect 1306 923 1325 926
rect 1346 923 1349 936
rect 1434 933 1437 996
rect 1450 936 1453 996
rect 1450 933 1469 936
rect 1514 933 1517 1016
rect 1530 933 1533 986
rect 1322 913 1325 923
rect 1306 796 1309 806
rect 1314 803 1317 826
rect 1338 813 1341 826
rect 1354 813 1357 926
rect 1410 873 1413 926
rect 1378 813 1381 856
rect 1450 853 1453 926
rect 1466 856 1469 933
rect 1458 853 1469 856
rect 1458 833 1461 853
rect 1386 813 1389 826
rect 1418 806 1421 816
rect 1306 793 1317 796
rect 1362 733 1365 746
rect 1226 723 1237 726
rect 1210 693 1221 696
rect 1210 636 1213 693
rect 1210 633 1221 636
rect 1218 613 1221 633
rect 1162 533 1189 536
rect 1018 363 1037 366
rect 1026 333 1029 346
rect 1034 333 1037 363
rect 1026 223 1029 326
rect 1042 323 1045 386
rect 1066 343 1069 406
rect 1106 403 1117 406
rect 1114 353 1117 403
rect 1050 263 1053 336
rect 1138 333 1141 416
rect 1146 413 1149 526
rect 1154 523 1165 526
rect 1194 523 1197 546
rect 1234 533 1237 723
rect 1242 703 1245 726
rect 1258 713 1261 726
rect 1338 706 1341 726
rect 1330 703 1341 706
rect 1346 723 1365 726
rect 1330 626 1333 703
rect 1250 533 1253 626
rect 1330 623 1341 626
rect 1346 623 1349 723
rect 1362 703 1373 706
rect 1394 703 1397 716
rect 1338 606 1341 623
rect 1362 613 1365 676
rect 1410 613 1413 806
rect 1418 803 1429 806
rect 1474 803 1485 806
rect 1426 786 1429 803
rect 1426 783 1437 786
rect 1474 783 1477 796
rect 1434 733 1437 783
rect 1490 736 1493 926
rect 1514 826 1517 926
rect 1514 823 1525 826
rect 1418 713 1421 726
rect 1442 716 1445 736
rect 1482 733 1493 736
rect 1434 673 1437 716
rect 1442 713 1453 716
rect 1482 713 1485 733
rect 1514 726 1517 816
rect 1522 805 1525 823
rect 1538 803 1541 1016
rect 1578 1013 1581 1026
rect 1586 1003 1589 1036
rect 1674 1023 1677 1066
rect 1686 1016 1689 1073
rect 1682 1013 1689 1016
rect 1546 923 1549 936
rect 1634 933 1637 946
rect 1586 813 1589 876
rect 1642 846 1645 936
rect 1650 883 1653 1006
rect 1658 866 1661 926
rect 1618 826 1621 846
rect 1634 843 1645 846
rect 1654 863 1661 866
rect 1634 826 1637 843
rect 1610 823 1621 826
rect 1630 823 1637 826
rect 1642 823 1645 836
rect 1490 723 1517 726
rect 1530 723 1533 736
rect 1450 656 1453 713
rect 1498 703 1501 716
rect 1506 703 1509 716
rect 1514 673 1517 716
rect 1442 653 1453 656
rect 1442 633 1445 653
rect 1330 603 1349 606
rect 1386 553 1389 606
rect 1250 506 1253 526
rect 1242 503 1253 506
rect 1242 436 1245 503
rect 1242 433 1253 436
rect 1170 423 1181 426
rect 1154 413 1173 416
rect 898 123 901 166
rect 946 123 949 206
rect 986 133 989 216
rect 1082 213 1085 326
rect 1170 323 1173 406
rect 1178 373 1181 423
rect 1250 413 1253 433
rect 1266 413 1269 526
rect 1314 523 1317 546
rect 1402 523 1405 596
rect 1498 586 1501 596
rect 1506 593 1509 606
rect 1514 586 1517 606
rect 1498 583 1517 586
rect 1410 523 1413 536
rect 1418 496 1421 526
rect 1410 493 1421 496
rect 1410 426 1413 493
rect 1410 423 1421 426
rect 1218 306 1221 396
rect 1210 303 1221 306
rect 1210 256 1213 303
rect 1226 263 1229 336
rect 1298 333 1301 406
rect 1210 253 1221 256
rect 1002 133 1005 166
rect 1042 163 1045 206
rect 1066 156 1069 206
rect 954 123 965 126
rect 1026 123 1029 136
rect 1042 123 1045 146
rect 1050 133 1053 156
rect 1066 153 1077 156
rect 1074 126 1077 153
rect 1082 133 1085 186
rect 1114 183 1117 206
rect 1122 163 1125 216
rect 1090 133 1093 146
rect 1138 133 1141 156
rect 1178 133 1181 226
rect 1218 223 1221 253
rect 1234 183 1237 216
rect 1242 203 1253 206
rect 1250 133 1253 203
rect 1266 196 1269 216
rect 1274 203 1277 226
rect 1282 213 1285 326
rect 1306 323 1309 376
rect 1354 333 1357 396
rect 1362 393 1365 406
rect 1394 333 1397 346
rect 1322 313 1325 326
rect 1330 213 1333 226
rect 1282 196 1285 206
rect 1266 193 1285 196
rect 1258 133 1261 156
rect 1266 143 1269 193
rect 1338 173 1341 216
rect 1386 213 1397 216
rect 1418 213 1421 423
rect 1426 413 1429 566
rect 1434 406 1437 416
rect 1426 403 1437 406
rect 1426 353 1429 403
rect 1442 376 1445 536
rect 1434 373 1445 376
rect 1434 343 1437 373
rect 1450 366 1453 406
rect 1466 403 1469 526
rect 1490 523 1493 536
rect 1530 533 1533 556
rect 1474 423 1477 436
rect 1442 363 1453 366
rect 1442 323 1445 363
rect 1474 306 1477 326
rect 1466 303 1477 306
rect 1466 246 1469 303
rect 1466 243 1477 246
rect 1074 123 1093 126
rect 1226 103 1229 126
rect 1354 113 1357 126
rect 1370 103 1373 136
rect 1402 133 1421 136
rect 1410 103 1413 126
rect 786 0 789 96
rect 1418 0 1421 133
rect 1426 123 1429 206
rect 1474 203 1477 243
rect 1482 223 1485 326
rect 1490 313 1493 516
rect 1514 413 1517 436
rect 1530 416 1533 526
rect 1530 413 1541 416
rect 1554 413 1557 806
rect 1610 756 1613 823
rect 1610 753 1621 756
rect 1618 733 1621 753
rect 1630 746 1633 823
rect 1630 743 1637 746
rect 1626 713 1629 726
rect 1634 696 1637 743
rect 1626 693 1637 696
rect 1626 626 1629 693
rect 1642 683 1645 806
rect 1654 796 1657 863
rect 1650 793 1657 796
rect 1626 623 1637 626
rect 1634 606 1637 623
rect 1578 533 1589 536
rect 1626 533 1629 606
rect 1634 603 1641 606
rect 1638 546 1641 603
rect 1634 543 1641 546
rect 1594 513 1597 526
rect 1634 523 1637 543
rect 1650 523 1653 793
rect 1666 733 1669 936
rect 1682 933 1685 1013
rect 1698 996 1701 1156
rect 1714 1133 1717 1183
rect 1734 1176 1737 1223
rect 1754 1206 1757 1296
rect 1762 1213 1765 1326
rect 1786 1323 1789 1336
rect 1794 1333 1797 1406
rect 1818 1403 1829 1406
rect 1834 1403 1837 1436
rect 1874 1433 1885 1436
rect 1842 1403 1845 1426
rect 1882 1413 1885 1433
rect 1778 1223 1781 1306
rect 1730 1173 1737 1176
rect 1722 1133 1725 1156
rect 1730 1136 1733 1173
rect 1746 1156 1749 1206
rect 1754 1203 1765 1206
rect 1802 1173 1805 1356
rect 1818 1323 1821 1403
rect 1898 1393 1901 1456
rect 1922 1446 1925 1523
rect 1938 1453 1941 1516
rect 1954 1486 1957 1526
rect 1970 1503 1973 1583
rect 1994 1536 1997 1556
rect 1986 1526 1989 1536
rect 1994 1533 2005 1536
rect 2018 1533 2021 1616
rect 2122 1613 2125 1726
rect 1978 1523 1997 1526
rect 2002 1523 2005 1533
rect 1954 1483 1965 1486
rect 1922 1443 1933 1446
rect 1914 1346 1917 1396
rect 1826 1233 1829 1336
rect 1834 1333 1837 1346
rect 1906 1343 1917 1346
rect 1810 1223 1837 1226
rect 1810 1213 1813 1223
rect 1818 1213 1829 1216
rect 1842 1213 1845 1316
rect 1882 1313 1885 1326
rect 1906 1303 1909 1343
rect 1738 1146 1741 1156
rect 1746 1153 1765 1156
rect 1738 1143 1749 1146
rect 1730 1133 1749 1136
rect 1714 1013 1717 1036
rect 1730 1033 1733 1056
rect 1738 1033 1741 1126
rect 1762 1123 1765 1153
rect 1810 1136 1813 1206
rect 1858 1205 1861 1216
rect 1802 1133 1813 1136
rect 1802 1056 1805 1133
rect 1802 1053 1813 1056
rect 1738 1013 1741 1026
rect 1698 993 1709 996
rect 1674 833 1677 926
rect 1690 923 1693 936
rect 1682 766 1685 886
rect 1706 836 1709 993
rect 1746 946 1749 1036
rect 1786 1013 1789 1036
rect 1674 763 1685 766
rect 1698 833 1709 836
rect 1730 943 1749 946
rect 1730 836 1733 943
rect 1754 846 1757 936
rect 1786 876 1789 916
rect 1794 906 1797 1026
rect 1810 1016 1813 1053
rect 1810 1013 1821 1016
rect 1826 1013 1829 1126
rect 1842 1053 1845 1146
rect 1850 1133 1853 1176
rect 1882 1133 1885 1216
rect 1930 1213 1933 1443
rect 1962 1356 1965 1483
rect 1986 1453 1989 1516
rect 2026 1466 2029 1516
rect 2034 1496 2037 1526
rect 2042 1516 2045 1536
rect 2050 1523 2053 1536
rect 2082 1533 2085 1596
rect 2106 1593 2109 1606
rect 2058 1516 2061 1526
rect 2042 1513 2061 1516
rect 2034 1493 2045 1496
rect 2018 1463 2029 1466
rect 1978 1403 1981 1416
rect 1954 1353 1965 1356
rect 1938 1196 1941 1306
rect 1954 1296 1957 1353
rect 1962 1333 1965 1346
rect 2010 1333 2013 1416
rect 1954 1293 1965 1296
rect 1962 1226 1965 1293
rect 1954 1223 1965 1226
rect 1954 1203 1957 1223
rect 1986 1213 1989 1326
rect 2018 1316 2021 1463
rect 2026 1413 2029 1456
rect 2042 1426 2045 1493
rect 2034 1423 2045 1426
rect 2034 1403 2037 1423
rect 2050 1403 2061 1406
rect 2026 1323 2029 1396
rect 2066 1393 2069 1426
rect 2034 1333 2037 1346
rect 2042 1343 2045 1366
rect 2138 1323 2141 1596
rect 2018 1313 2037 1316
rect 2034 1293 2037 1313
rect 2058 1226 2061 1296
rect 2058 1223 2069 1226
rect 1970 1203 1997 1206
rect 1938 1193 1949 1196
rect 2042 1193 2045 1206
rect 1938 1186 1941 1193
rect 1922 1183 1941 1186
rect 1922 1133 1925 1183
rect 1946 1166 1949 1186
rect 1942 1163 1949 1166
rect 1858 1123 1877 1126
rect 1906 1103 1909 1116
rect 1930 1086 1933 1126
rect 1922 1083 1933 1086
rect 1942 1086 1945 1163
rect 2010 1133 2013 1186
rect 2026 1133 2029 1186
rect 2050 1183 2053 1216
rect 2066 1176 2069 1223
rect 2058 1173 2069 1176
rect 1986 1113 1989 1126
rect 2026 1103 2029 1126
rect 1942 1083 1949 1086
rect 1810 976 1813 1006
rect 1802 973 1813 976
rect 1802 913 1805 973
rect 1818 966 1821 1013
rect 1810 963 1821 966
rect 1810 923 1813 963
rect 1834 936 1837 1036
rect 1842 996 1845 1026
rect 1842 993 1853 996
rect 1818 933 1837 936
rect 1850 926 1853 993
rect 1922 976 1925 1083
rect 1946 1003 1949 1083
rect 1922 973 1933 976
rect 1930 956 1933 973
rect 1930 953 1949 956
rect 1818 906 1821 926
rect 1794 903 1821 906
rect 1786 873 1797 876
rect 1778 846 1781 866
rect 1754 843 1765 846
rect 1730 833 1749 836
rect 1674 623 1677 763
rect 1698 746 1701 833
rect 1714 813 1741 816
rect 1682 723 1685 746
rect 1690 743 1701 746
rect 1690 706 1693 743
rect 1698 716 1701 736
rect 1706 723 1709 766
rect 1730 736 1733 806
rect 1746 803 1749 833
rect 1762 796 1765 843
rect 1754 793 1765 796
rect 1774 843 1781 846
rect 1774 796 1777 843
rect 1794 826 1797 873
rect 1786 823 1797 826
rect 1818 823 1821 903
rect 1842 923 1853 926
rect 1906 923 1909 936
rect 1786 803 1789 823
rect 1842 816 1845 923
rect 1774 793 1781 796
rect 1802 793 1805 806
rect 1714 716 1717 736
rect 1698 713 1717 716
rect 1722 733 1733 736
rect 1690 703 1701 706
rect 1610 503 1613 516
rect 1650 413 1653 516
rect 1666 503 1669 526
rect 1506 393 1509 406
rect 1514 403 1525 406
rect 1530 326 1533 406
rect 1538 386 1541 413
rect 1538 383 1549 386
rect 1514 323 1533 326
rect 1514 256 1517 323
rect 1506 253 1517 256
rect 1506 213 1509 253
rect 1482 186 1485 206
rect 1466 183 1485 186
rect 1434 113 1437 126
rect 1466 123 1469 183
rect 1474 133 1477 156
rect 1530 153 1533 206
rect 1482 123 1485 136
rect 1546 133 1549 383
rect 1562 333 1565 346
rect 1586 343 1589 406
rect 1602 326 1605 406
rect 1674 346 1677 526
rect 1682 513 1685 526
rect 1690 496 1693 696
rect 1686 493 1693 496
rect 1686 426 1689 493
rect 1686 423 1693 426
rect 1698 423 1701 703
rect 1706 656 1709 713
rect 1722 676 1725 733
rect 1730 713 1733 726
rect 1738 693 1741 746
rect 1754 743 1757 793
rect 1722 673 1733 676
rect 1706 653 1717 656
rect 1714 576 1717 653
rect 1706 573 1717 576
rect 1706 496 1709 573
rect 1730 556 1733 673
rect 1762 603 1765 616
rect 1778 605 1781 793
rect 1810 676 1813 736
rect 1818 713 1821 816
rect 1842 813 1853 816
rect 1842 753 1845 806
rect 1826 723 1829 736
rect 1834 733 1837 746
rect 1810 673 1821 676
rect 1730 553 1741 556
rect 1714 503 1717 546
rect 1706 493 1717 496
rect 1682 393 1685 406
rect 1690 403 1693 423
rect 1666 343 1677 346
rect 1666 333 1669 343
rect 1682 336 1685 366
rect 1674 333 1685 336
rect 1586 323 1605 326
rect 1586 213 1589 323
rect 1546 113 1549 126
rect 1554 103 1557 126
rect 1562 116 1565 206
rect 1562 113 1573 116
rect 1578 113 1581 126
rect 1594 123 1597 156
rect 1610 113 1613 206
rect 1618 203 1621 256
rect 1666 133 1669 246
rect 1698 113 1701 416
rect 1706 396 1709 426
rect 1714 423 1717 493
rect 1738 436 1741 553
rect 1778 493 1781 526
rect 1722 433 1741 436
rect 1722 413 1725 433
rect 1786 423 1789 526
rect 1802 456 1805 616
rect 1818 516 1821 673
rect 1850 626 1853 813
rect 1898 793 1901 886
rect 1930 883 1933 936
rect 1922 776 1925 816
rect 1946 813 1949 953
rect 1954 943 1957 966
rect 1970 946 1973 1016
rect 1962 943 1973 946
rect 1962 936 1965 943
rect 1954 933 1965 936
rect 1978 933 1981 956
rect 1986 943 1989 1076
rect 2026 1003 2029 1016
rect 2034 1003 2037 1116
rect 2058 1113 2061 1173
rect 1954 923 1957 933
rect 1978 826 1981 926
rect 1978 823 1989 826
rect 1986 803 1989 823
rect 1994 793 1997 936
rect 2010 923 2013 966
rect 2034 963 2037 996
rect 2026 863 2029 936
rect 2050 923 2053 1006
rect 2066 933 2069 986
rect 2114 933 2117 1006
rect 2138 933 2141 956
rect 2146 923 2149 976
rect 2010 803 2013 816
rect 2018 813 2021 826
rect 1906 773 1925 776
rect 1858 703 1861 726
rect 1866 723 1869 746
rect 1898 723 1901 736
rect 1906 733 1909 773
rect 1898 636 1901 716
rect 1914 713 1917 726
rect 1922 723 1925 756
rect 2002 733 2005 796
rect 2026 763 2029 816
rect 2058 813 2061 826
rect 1846 623 1853 626
rect 1882 633 1901 636
rect 1846 536 1849 623
rect 1846 533 1853 536
rect 1858 533 1861 616
rect 1882 546 1885 633
rect 1914 605 1917 616
rect 1938 613 1941 726
rect 1954 713 1957 726
rect 2026 686 2029 736
rect 2050 723 2053 806
rect 2066 713 2069 826
rect 2114 806 2117 916
rect 2114 803 2125 806
rect 2106 703 2109 766
rect 2130 736 2133 746
rect 2114 733 2133 736
rect 2114 723 2117 733
rect 2026 683 2037 686
rect 1882 543 1901 546
rect 1810 513 1829 516
rect 1850 513 1853 533
rect 1794 453 1805 456
rect 1738 403 1741 416
rect 1706 393 1717 396
rect 1714 336 1717 393
rect 1754 383 1757 406
rect 1706 333 1717 336
rect 1706 313 1709 333
rect 1770 323 1773 346
rect 1786 333 1789 406
rect 1794 403 1797 453
rect 1818 413 1821 506
rect 1874 423 1877 526
rect 1898 523 1901 543
rect 1914 533 1917 556
rect 1954 536 1957 606
rect 1930 533 1957 536
rect 1834 383 1837 406
rect 1786 216 1789 326
rect 1842 306 1845 406
rect 1858 366 1861 386
rect 1834 303 1845 306
rect 1854 363 1861 366
rect 1834 246 1837 303
rect 1854 286 1857 363
rect 1882 323 1885 406
rect 1898 393 1901 416
rect 1906 383 1909 526
rect 1930 523 1933 533
rect 1946 503 1949 516
rect 1954 423 1957 526
rect 1962 523 1965 546
rect 1970 503 1973 526
rect 1978 513 1981 526
rect 1986 506 1989 616
rect 1994 553 1997 636
rect 2034 605 2037 683
rect 2114 666 2117 716
rect 2122 713 2125 726
rect 2098 663 2117 666
rect 1978 503 1989 506
rect 1854 283 1861 286
rect 1834 243 1845 246
rect 1802 223 1805 236
rect 1810 223 1837 226
rect 1706 206 1709 216
rect 1706 203 1725 206
rect 1570 0 1573 113
rect 1730 3 1733 216
rect 1786 213 1793 216
rect 1810 213 1813 223
rect 1762 133 1765 196
rect 1770 106 1773 126
rect 1762 103 1773 106
rect 1762 16 1765 103
rect 1778 83 1781 206
rect 1790 76 1793 213
rect 1810 183 1813 206
rect 1818 203 1821 216
rect 1842 213 1845 243
rect 1834 123 1837 206
rect 1850 193 1853 216
rect 1858 183 1861 283
rect 1874 196 1877 216
rect 1874 193 1885 196
rect 1858 133 1861 146
rect 1882 106 1885 193
rect 1874 103 1885 106
rect 1786 73 1793 76
rect 1762 13 1773 16
rect 1714 0 1733 3
rect 1770 0 1773 13
rect 1786 0 1789 73
rect 1802 0 1805 86
rect 1850 0 1853 86
rect 1874 83 1877 103
rect 1906 83 1909 196
rect 1922 143 1925 356
rect 1978 353 1981 503
rect 2002 483 2005 516
rect 2018 473 2021 536
rect 2026 513 2029 536
rect 2034 526 2037 576
rect 2058 533 2061 616
rect 2098 576 2101 663
rect 2090 573 2101 576
rect 2034 523 2053 526
rect 2066 503 2069 516
rect 2082 513 2085 526
rect 2002 413 2005 426
rect 2058 413 2061 476
rect 2066 376 2069 426
rect 2090 423 2093 573
rect 2114 533 2117 616
rect 2122 613 2125 706
rect 2146 613 2149 626
rect 2098 503 2101 526
rect 2062 373 2069 376
rect 1970 313 1973 326
rect 1970 223 1973 236
rect 1978 213 1981 346
rect 1994 333 1997 356
rect 2042 323 2045 346
rect 2062 316 2065 373
rect 2074 323 2077 366
rect 2082 333 2085 386
rect 2090 323 2093 406
rect 2098 326 2101 416
rect 2106 363 2109 406
rect 2106 333 2109 346
rect 2114 333 2117 356
rect 2098 323 2109 326
rect 2062 313 2069 316
rect 2106 313 2109 323
rect 2066 233 2069 313
rect 2130 303 2133 326
rect 2098 223 2101 236
rect 1946 123 1949 206
rect 1954 193 1957 206
rect 1970 183 1973 206
rect 1986 133 1989 146
rect 2042 133 2045 146
rect 2074 123 2077 206
rect 2082 163 2085 206
rect 2122 123 2125 166
rect 1930 0 1933 86
rect 2160 37 2180 2003
rect 2184 13 2204 2027
<< metal3 >>
rect 977 1972 1070 1977
rect 513 1962 574 1967
rect 1217 1962 1262 1967
rect 625 1952 734 1957
rect 1049 1952 1118 1957
rect 113 1942 230 1947
rect 265 1942 366 1947
rect 537 1942 622 1947
rect 777 1942 822 1947
rect 953 1942 1006 1947
rect 1105 1932 1142 1937
rect 193 1922 222 1927
rect 217 1917 222 1922
rect 297 1922 526 1927
rect 297 1917 302 1922
rect 217 1912 302 1917
rect 521 1917 526 1922
rect 633 1922 918 1927
rect 1041 1922 1134 1927
rect 1153 1922 1158 1957
rect 1417 1952 1494 1957
rect 1665 1952 1726 1957
rect 1417 1947 1422 1952
rect 1233 1942 1278 1947
rect 1377 1942 1422 1947
rect 1489 1947 1494 1952
rect 1489 1942 1518 1947
rect 1553 1942 1662 1947
rect 1809 1942 1934 1947
rect 1977 1942 2062 1947
rect 1865 1932 1894 1937
rect 1889 1927 1894 1932
rect 2001 1932 2030 1937
rect 2001 1927 2006 1932
rect 1433 1922 1494 1927
rect 1585 1922 1678 1927
rect 1889 1922 2006 1927
rect 633 1917 638 1922
rect 521 1912 638 1917
rect 1137 1912 1342 1917
rect 1497 1902 1582 1907
rect 1209 1897 1310 1902
rect 1185 1892 1214 1897
rect 1305 1892 1334 1897
rect 1201 1882 1230 1887
rect 1225 1877 1230 1882
rect 1345 1882 1510 1887
rect 1345 1877 1350 1882
rect 1225 1872 1350 1877
rect 1505 1877 1510 1882
rect 1593 1882 1830 1887
rect 1881 1882 1942 1887
rect 1985 1882 2014 1887
rect 1593 1877 1598 1882
rect 1505 1872 1598 1877
rect 1721 1872 1766 1877
rect 921 1862 1022 1867
rect 1249 1852 1286 1857
rect 881 1832 918 1837
rect 1153 1832 1206 1837
rect 177 1822 302 1827
rect 369 1822 414 1827
rect 961 1822 1006 1827
rect 1177 1822 1238 1827
rect 1257 1822 1350 1827
rect 2033 1822 2062 1827
rect 1257 1817 1262 1822
rect 569 1812 654 1817
rect 977 1807 982 1817
rect 1145 1812 1262 1817
rect 1345 1817 1350 1822
rect 1345 1812 1374 1817
rect 1681 1812 1734 1817
rect 1777 1812 2046 1817
rect 697 1802 878 1807
rect 937 1802 982 1807
rect 1025 1802 1118 1807
rect 1225 1802 1550 1807
rect 1025 1797 1030 1802
rect 193 1792 366 1797
rect 377 1792 446 1797
rect 521 1792 566 1797
rect 633 1792 670 1797
rect 777 1792 894 1797
rect 905 1792 1030 1797
rect 1113 1797 1118 1802
rect 1113 1792 1422 1797
rect 81 1782 198 1787
rect 217 1782 270 1787
rect 353 1782 390 1787
rect 953 1782 982 1787
rect 977 1777 982 1782
rect 1041 1782 1158 1787
rect 1209 1782 1262 1787
rect 1561 1782 1614 1787
rect 1041 1777 1046 1782
rect 977 1772 1046 1777
rect 193 1762 230 1767
rect 1393 1762 1430 1767
rect 361 1742 590 1747
rect 321 1732 350 1737
rect 345 1727 350 1732
rect 457 1732 486 1737
rect 457 1727 462 1732
rect 345 1722 462 1727
rect 553 1722 582 1727
rect 713 1722 758 1727
rect 209 1712 278 1717
rect 769 1712 774 1757
rect 945 1752 1022 1757
rect 945 1747 950 1752
rect 825 1742 950 1747
rect 1017 1747 1022 1752
rect 1065 1752 1222 1757
rect 1649 1752 1678 1757
rect 1969 1752 1990 1757
rect 1065 1747 1070 1752
rect 1017 1742 1070 1747
rect 1217 1747 1222 1752
rect 1217 1742 1246 1747
rect 961 1732 990 1737
rect 985 1727 990 1732
rect 1097 1732 1150 1737
rect 1193 1732 1286 1737
rect 1729 1732 1894 1737
rect 1097 1727 1102 1732
rect 985 1722 1102 1727
rect 1585 1722 1726 1727
rect 2041 1722 2126 1727
rect 1121 1712 1206 1717
rect 1929 1712 2038 1717
rect 281 1702 350 1707
rect 433 1702 486 1707
rect 649 1702 702 1707
rect 697 1697 702 1702
rect 769 1702 814 1707
rect 769 1697 774 1702
rect 697 1692 774 1697
rect 793 1692 902 1697
rect 1433 1662 1614 1667
rect 737 1652 814 1657
rect 1017 1652 1054 1657
rect 737 1647 742 1652
rect 617 1642 742 1647
rect 809 1647 814 1652
rect 1433 1647 1438 1662
rect 809 1642 838 1647
rect 1313 1642 1390 1647
rect 1409 1642 1438 1647
rect 1609 1647 1614 1662
rect 1609 1642 1806 1647
rect 1313 1637 1318 1642
rect 145 1632 542 1637
rect 625 1632 654 1637
rect 1025 1632 1046 1637
rect 1289 1632 1318 1637
rect 1385 1637 1390 1642
rect 1385 1632 1598 1637
rect 233 1622 270 1627
rect 753 1622 862 1627
rect 537 1612 662 1617
rect 945 1612 998 1617
rect 585 1602 646 1607
rect 649 1592 822 1597
rect 849 1592 894 1597
rect 921 1582 958 1587
rect 1041 1582 1046 1632
rect 1073 1622 1230 1627
rect 1281 1622 1382 1627
rect 1249 1612 1270 1617
rect 1417 1612 1510 1617
rect 1553 1612 1622 1617
rect 1249 1592 1478 1597
rect 1537 1592 1774 1597
rect 1817 1592 1982 1597
rect 2105 1592 2142 1597
rect 1529 1582 1598 1587
rect 441 1572 502 1577
rect 1217 1572 1326 1577
rect 481 1562 526 1567
rect 1761 1562 1838 1567
rect 1761 1557 1766 1562
rect 1689 1552 1766 1557
rect 1833 1557 1838 1562
rect 1833 1552 1998 1557
rect 81 1542 438 1547
rect 449 1542 510 1547
rect 985 1542 1030 1547
rect 1073 1542 1142 1547
rect 1225 1542 1334 1547
rect 1225 1537 1230 1542
rect 841 1532 974 1537
rect 969 1527 974 1532
rect 1105 1532 1230 1537
rect 1329 1537 1334 1542
rect 1441 1542 1526 1547
rect 1593 1542 1822 1547
rect 1441 1537 1446 1542
rect 1329 1532 1446 1537
rect 1521 1537 1526 1542
rect 1521 1532 1582 1537
rect 1105 1527 1110 1532
rect 529 1522 566 1527
rect 969 1522 1110 1527
rect 1265 1522 1318 1527
rect 1457 1522 1502 1527
rect 1577 1517 1582 1532
rect 1705 1532 1750 1537
rect 1985 1532 2054 1537
rect 1705 1517 1710 1532
rect 1729 1522 1734 1532
rect 2001 1522 2038 1527
rect 497 1512 526 1517
rect 1241 1512 1278 1517
rect 1481 1512 1510 1517
rect 1577 1512 1710 1517
rect 1809 1512 1854 1517
rect 177 1502 350 1507
rect 441 1502 486 1507
rect 481 1497 486 1502
rect 577 1502 774 1507
rect 1129 1502 1326 1507
rect 1801 1502 2030 1507
rect 577 1497 582 1502
rect 481 1492 582 1497
rect 897 1492 1118 1497
rect 1113 1477 1118 1492
rect 1273 1492 1366 1497
rect 1273 1477 1278 1492
rect 1817 1482 1902 1487
rect 1113 1472 1278 1477
rect 1897 1452 1942 1457
rect 1985 1452 2030 1457
rect 937 1442 1086 1447
rect 241 1432 430 1437
rect 481 1432 662 1437
rect 1025 1432 1382 1437
rect 1809 1432 1838 1437
rect 233 1422 262 1427
rect 713 1422 814 1427
rect 1489 1422 1534 1427
rect 1649 1422 1734 1427
rect 1801 1422 1846 1427
rect 2001 1422 2220 1427
rect 713 1417 718 1422
rect 193 1412 230 1417
rect 377 1412 414 1417
rect 449 1412 582 1417
rect 577 1407 582 1412
rect 673 1412 718 1417
rect 809 1417 814 1422
rect 1649 1417 1654 1422
rect 1729 1417 1734 1422
rect 2001 1417 2006 1422
rect 809 1412 886 1417
rect 1009 1412 1030 1417
rect 1473 1412 1654 1417
rect 1689 1412 1718 1417
rect 1729 1412 2006 1417
rect 673 1407 678 1412
rect 577 1402 678 1407
rect 1977 1402 2054 1407
rect 129 1392 222 1397
rect 729 1392 862 1397
rect 905 1392 974 1397
rect 1649 1392 1686 1397
rect 2025 1392 2070 1397
rect 385 1382 422 1387
rect 705 1382 830 1387
rect 977 1382 1094 1387
rect 193 1372 254 1377
rect 473 1372 550 1377
rect 473 1367 478 1372
rect 425 1362 478 1367
rect 545 1367 550 1372
rect 545 1362 574 1367
rect 1209 1362 1294 1367
rect 1313 1362 1430 1367
rect 1465 1362 1502 1367
rect 2009 1362 2046 1367
rect 1313 1357 1318 1362
rect 489 1342 550 1347
rect 689 1342 782 1347
rect 161 1332 278 1337
rect 321 1322 374 1327
rect 393 1322 478 1327
rect 321 1317 326 1322
rect 473 1317 478 1322
rect 553 1322 590 1327
rect 801 1322 806 1357
rect 1137 1352 1318 1357
rect 1425 1357 1430 1362
rect 1425 1352 1542 1357
rect 1673 1352 1806 1357
rect 945 1342 966 1347
rect 1225 1342 1254 1347
rect 1329 1342 1438 1347
rect 1249 1337 1334 1342
rect 1433 1337 1438 1342
rect 1529 1342 1582 1347
rect 1777 1342 1838 1347
rect 1961 1342 2038 1347
rect 1529 1337 1534 1342
rect 1129 1332 1166 1337
rect 1433 1332 1534 1337
rect 1793 1332 1830 1337
rect 897 1322 958 1327
rect 1049 1322 1118 1327
rect 1249 1322 1270 1327
rect 1361 1322 1398 1327
rect 1553 1322 1614 1327
rect 1705 1322 1790 1327
rect 1985 1322 1990 1342
rect 553 1317 558 1322
rect 1393 1317 1398 1322
rect 177 1312 326 1317
rect 337 1292 342 1317
rect 473 1312 558 1317
rect 577 1312 622 1317
rect 753 1312 1070 1317
rect 1393 1312 1510 1317
rect 1841 1312 1886 1317
rect 369 1302 422 1307
rect 641 1302 710 1307
rect 1025 1302 1286 1307
rect 1377 1302 1406 1307
rect 1401 1297 1406 1302
rect 1473 1302 1574 1307
rect 1721 1302 1862 1307
rect 1905 1302 1942 1307
rect 1473 1297 1478 1302
rect 1857 1297 1862 1302
rect 1065 1292 1174 1297
rect 1169 1287 1174 1292
rect 1233 1292 1286 1297
rect 1401 1292 1478 1297
rect 1577 1292 1758 1297
rect 1857 1292 1878 1297
rect 1233 1287 1238 1292
rect 73 1282 278 1287
rect 569 1282 678 1287
rect 1097 1282 1150 1287
rect 1169 1282 1238 1287
rect 73 1267 78 1282
rect 0 1262 78 1267
rect 273 1267 278 1282
rect 1281 1277 1286 1292
rect 1577 1277 1582 1292
rect 1873 1287 1878 1292
rect 1953 1292 2062 1297
rect 1953 1287 1958 1292
rect 1873 1282 1958 1287
rect 1281 1272 1582 1277
rect 1601 1272 1630 1277
rect 1625 1267 1630 1272
rect 1769 1272 1846 1277
rect 1769 1267 1774 1272
rect 273 1262 838 1267
rect 1625 1262 1774 1267
rect 1841 1267 1846 1272
rect 2073 1272 2220 1277
rect 2073 1267 2078 1272
rect 1841 1262 2078 1267
rect 89 1252 262 1257
rect 1313 1242 1342 1247
rect 209 1232 254 1237
rect 729 1232 790 1237
rect 265 1222 318 1227
rect 753 1222 822 1227
rect 225 1212 294 1217
rect 417 1212 446 1217
rect 1329 1212 1374 1217
rect 1825 1212 1830 1237
rect 1857 1212 1934 1217
rect 1105 1202 1150 1207
rect 1649 1202 1686 1207
rect 1761 1202 1814 1207
rect 673 1192 926 1197
rect 1137 1192 1198 1197
rect 1449 1192 1638 1197
rect 1633 1187 1638 1192
rect 1697 1192 1814 1197
rect 1937 1192 2046 1197
rect 1697 1187 1702 1192
rect 793 1182 846 1187
rect 1633 1182 1702 1187
rect 1809 1187 1814 1192
rect 1809 1182 2014 1187
rect 2025 1182 2054 1187
rect 1169 1172 1342 1177
rect 1801 1172 1854 1177
rect 785 1162 894 1167
rect 1169 1162 1334 1167
rect 1345 1162 1366 1167
rect 785 1157 790 1162
rect 137 1152 214 1157
rect 489 1152 566 1157
rect 657 1152 790 1157
rect 889 1157 894 1162
rect 889 1152 1158 1157
rect 1153 1147 1158 1152
rect 1289 1152 1742 1157
rect 1289 1147 1294 1152
rect 233 1142 262 1147
rect 401 1142 550 1147
rect 281 1132 382 1137
rect 201 1127 286 1132
rect 377 1127 462 1132
rect 0 1122 206 1127
rect 457 1122 542 1127
rect 217 1112 358 1117
rect 409 1112 446 1117
rect 625 1112 750 1117
rect 801 1112 806 1147
rect 841 1142 878 1147
rect 1153 1142 1294 1147
rect 1033 1122 1110 1127
rect 1313 1122 1318 1147
rect 1761 1142 1846 1147
rect 1865 1132 2054 1137
rect 1865 1127 1870 1132
rect 1337 1122 1422 1127
rect 1337 1117 1342 1122
rect 1289 1112 1342 1117
rect 1417 1117 1422 1122
rect 1841 1122 1870 1127
rect 2049 1127 2054 1132
rect 2049 1122 2220 1127
rect 1841 1117 1846 1122
rect 1417 1112 1846 1117
rect 1985 1112 2038 1117
rect 625 1107 630 1112
rect 233 1102 262 1107
rect 257 1097 262 1102
rect 393 1102 446 1107
rect 393 1097 398 1102
rect 257 1092 398 1097
rect 441 1097 446 1102
rect 553 1102 630 1107
rect 761 1102 782 1107
rect 1233 1102 1406 1107
rect 1905 1102 2030 1107
rect 553 1097 558 1102
rect 441 1092 558 1097
rect 1481 1082 1654 1087
rect 1161 1072 1262 1077
rect 1161 1067 1166 1072
rect 881 1062 1166 1067
rect 1257 1067 1262 1072
rect 1297 1072 1374 1077
rect 1297 1067 1302 1072
rect 1257 1062 1302 1067
rect 1369 1067 1374 1072
rect 1481 1067 1486 1082
rect 1369 1062 1486 1067
rect 1649 1067 1654 1082
rect 1985 1072 2220 1077
rect 1649 1062 1678 1067
rect 209 1052 462 1057
rect 1177 1052 1246 1057
rect 1497 1052 1638 1057
rect 1705 1052 1734 1057
rect 1841 1052 1990 1057
rect 209 1037 214 1052
rect 177 1032 214 1037
rect 457 1037 462 1052
rect 1633 1047 1710 1052
rect 1313 1042 1358 1047
rect 457 1032 486 1037
rect 945 1032 1102 1037
rect 1281 1032 1334 1037
rect 1505 1032 1590 1037
rect 1713 1032 1790 1037
rect 945 1027 950 1032
rect 225 1022 286 1027
rect 305 1022 446 1027
rect 537 1022 630 1027
rect 777 1022 910 1027
rect 921 1022 950 1027
rect 1097 1027 1102 1032
rect 1097 1022 1150 1027
rect 1305 1022 1462 1027
rect 1577 1022 1718 1027
rect 1737 1022 1830 1027
rect 457 1012 510 1017
rect 561 1012 766 1017
rect 913 1012 1142 1017
rect 761 1007 918 1012
rect 1713 1007 1718 1022
rect 1817 1012 1846 1017
rect 1817 1007 1822 1012
rect 433 1002 630 1007
rect 1113 1002 1214 1007
rect 1713 1002 1822 1007
rect 2025 1002 2054 1007
rect 241 992 318 997
rect 465 992 502 997
rect 745 992 774 997
rect 769 987 774 992
rect 881 992 910 997
rect 1017 992 1062 997
rect 881 987 886 992
rect 489 982 550 987
rect 769 982 886 987
rect 1057 987 1062 992
rect 1169 992 1438 997
rect 1937 992 2006 997
rect 1169 987 1174 992
rect 1937 987 1942 992
rect 1057 982 1174 987
rect 1529 982 1942 987
rect 2001 987 2006 992
rect 2001 982 2070 987
rect 2145 972 2220 977
rect 1953 962 1990 967
rect 2009 962 2038 967
rect 209 952 238 957
rect 441 952 558 957
rect 577 952 790 957
rect 1977 952 2220 957
rect 577 947 582 952
rect 121 942 182 947
rect 361 942 438 947
rect 457 942 582 947
rect 785 947 790 952
rect 785 942 1030 947
rect 1257 942 1318 947
rect 1369 942 1526 947
rect 1369 937 1374 942
rect 201 932 342 937
rect 737 932 774 937
rect 1345 932 1374 937
rect 1521 937 1526 942
rect 1521 932 1550 937
rect 1633 932 1694 937
rect 1905 932 2054 937
rect 2065 932 2220 937
rect 201 927 206 932
rect 0 922 206 927
rect 337 927 342 932
rect 337 922 686 927
rect 777 922 814 927
rect 1169 922 1294 927
rect 169 912 238 917
rect 297 912 326 917
rect 721 912 1062 917
rect 1257 912 1286 917
rect 1321 912 2220 917
rect 721 907 726 912
rect 153 902 182 907
rect 177 887 182 902
rect 337 902 422 907
rect 489 902 726 907
rect 1065 902 1182 907
rect 337 887 342 902
rect 1377 897 1494 902
rect 729 892 798 897
rect 1353 892 1382 897
rect 1489 892 1518 897
rect 1537 892 1606 897
rect 1537 887 1542 892
rect 177 882 342 887
rect 473 882 694 887
rect 1209 882 1542 887
rect 1601 887 1606 892
rect 1601 882 1686 887
rect 1897 882 2030 887
rect 2113 882 2220 887
rect 849 872 1118 877
rect 1409 872 1590 877
rect 849 857 854 872
rect 385 852 854 857
rect 1113 857 1118 872
rect 1137 862 1478 867
rect 1601 862 1782 867
rect 2025 862 2220 867
rect 1473 857 1606 862
rect 1113 852 1190 857
rect 1377 852 1454 857
rect 209 842 238 847
rect 793 842 1102 847
rect 1185 842 1214 847
rect 1289 842 1486 847
rect 1097 837 1190 842
rect 1481 837 1486 842
rect 1593 842 1622 847
rect 1993 842 2086 847
rect 1593 837 1598 842
rect 2081 837 2086 842
rect 2193 842 2220 847
rect 2193 837 2198 842
rect 185 832 230 837
rect 409 832 494 837
rect 785 832 854 837
rect 1441 832 1462 837
rect 1481 832 1598 837
rect 1641 832 1678 837
rect 2081 832 2198 837
rect 201 822 294 827
rect 585 822 654 827
rect 969 822 1158 827
rect 1193 822 1318 827
rect 1337 822 1390 827
rect 585 817 590 822
rect 0 812 590 817
rect 649 817 654 822
rect 1441 817 1446 832
rect 1873 822 1974 827
rect 2017 822 2062 827
rect 1873 817 1878 822
rect 649 812 686 817
rect 1417 812 1446 817
rect 1849 812 1878 817
rect 1969 817 1974 822
rect 1969 812 2014 817
rect 257 802 326 807
rect 601 802 638 807
rect 833 802 854 807
rect 961 802 998 807
rect 1409 802 1478 807
rect 153 792 214 797
rect 353 792 390 797
rect 1089 792 1310 797
rect 1801 792 1846 797
rect 1897 792 2006 797
rect 457 782 518 787
rect 1473 782 1670 787
rect 1825 772 1942 777
rect 1825 767 1830 772
rect 97 762 134 767
rect 545 762 662 767
rect 993 762 1078 767
rect 993 757 998 762
rect 121 752 158 757
rect 369 752 558 757
rect 969 752 998 757
rect 1073 757 1078 762
rect 1121 762 1342 767
rect 1705 762 1830 767
rect 1937 767 1942 772
rect 1937 762 2110 767
rect 1073 752 1102 757
rect 1121 747 1126 762
rect 169 742 238 747
rect 265 742 302 747
rect 361 742 406 747
rect 481 742 510 747
rect 849 742 966 747
rect 1089 742 1126 747
rect 1337 747 1342 762
rect 1401 752 1550 757
rect 1841 752 1926 757
rect 1337 742 1366 747
rect 1401 737 1406 752
rect 529 732 606 737
rect 785 732 886 737
rect 529 727 534 732
rect 417 722 534 727
rect 601 727 606 732
rect 881 727 886 732
rect 977 732 1078 737
rect 977 727 982 732
rect 601 722 630 727
rect 881 722 982 727
rect 1073 727 1078 732
rect 1137 732 1326 737
rect 1137 727 1142 732
rect 1073 722 1142 727
rect 1321 727 1326 732
rect 1385 732 1406 737
rect 1545 737 1550 752
rect 1681 742 1870 747
rect 2129 742 2220 747
rect 1545 732 1702 737
rect 1385 727 1390 732
rect 2049 727 2142 732
rect 1321 722 1390 727
rect 1417 722 1534 727
rect 1825 722 1854 727
rect 1897 722 1942 727
rect 1969 722 2054 727
rect 2137 722 2220 727
rect 417 717 422 722
rect 145 712 174 717
rect 281 712 422 717
rect 433 712 566 717
rect 641 712 710 717
rect 745 712 862 717
rect 1217 712 1262 717
rect 1481 712 1510 717
rect 1625 712 1822 717
rect 1913 712 1958 717
rect 561 707 646 712
rect 705 707 710 712
rect 1969 707 1974 722
rect 2065 712 2126 717
rect 705 702 774 707
rect 809 702 1366 707
rect 1393 702 1502 707
rect 1857 702 1974 707
rect 2105 702 2126 707
rect 609 692 638 697
rect 633 687 638 692
rect 697 692 806 697
rect 1689 692 1742 697
rect 697 687 702 692
rect 1345 687 1534 692
rect 633 682 702 687
rect 1113 682 1350 687
rect 1529 682 1646 687
rect 1361 672 1518 677
rect 721 662 806 667
rect 721 657 726 662
rect 129 652 302 657
rect 513 652 582 657
rect 697 652 726 657
rect 801 657 806 662
rect 801 652 1118 657
rect 1137 652 1270 657
rect 513 647 518 652
rect 465 642 518 647
rect 577 647 582 652
rect 577 642 614 647
rect 1137 637 1142 652
rect 737 632 790 637
rect 961 632 990 637
rect 985 627 990 632
rect 1105 632 1142 637
rect 1265 637 1270 652
rect 2129 642 2198 647
rect 2129 637 2134 642
rect 1265 632 1446 637
rect 1993 632 2134 637
rect 2193 637 2198 642
rect 2193 632 2220 637
rect 1105 627 1110 632
rect 153 622 182 627
rect 209 622 382 627
rect 401 622 430 627
rect 529 622 566 627
rect 841 622 894 627
rect 985 622 1110 627
rect 1129 622 1254 627
rect 1801 622 1894 627
rect 1801 617 1806 622
rect 441 612 686 617
rect 1777 612 1806 617
rect 1889 617 1894 622
rect 2145 617 2150 627
rect 1889 612 2038 617
rect 2145 612 2220 617
rect 1761 602 1958 607
rect 353 597 470 602
rect 81 592 118 597
rect 177 592 238 597
rect 265 592 358 597
rect 465 592 622 597
rect 1161 592 1382 597
rect 1401 592 1510 597
rect 1857 592 1886 597
rect 1969 592 2220 597
rect 385 582 454 587
rect 529 582 534 592
rect 1161 587 1166 592
rect 857 582 1166 587
rect 1377 587 1382 592
rect 1881 587 1974 592
rect 1377 582 1398 587
rect 1393 577 1398 582
rect 641 572 790 577
rect 1393 572 2038 577
rect 2113 572 2220 577
rect 641 567 646 572
rect 553 562 646 567
rect 553 557 558 562
rect 457 552 558 557
rect 785 557 790 572
rect 921 562 998 567
rect 1177 562 1430 567
rect 921 557 926 562
rect 785 552 926 557
rect 993 557 998 562
rect 993 552 1046 557
rect 1385 552 1534 557
rect 1913 552 1998 557
rect 1233 547 1366 552
rect 321 542 366 547
rect 561 542 654 547
rect 689 542 774 547
rect 937 542 1238 547
rect 1361 542 1718 547
rect 1961 542 2220 547
rect 769 537 854 542
rect 937 537 942 542
rect 849 532 942 537
rect 961 532 998 537
rect 1249 532 1414 537
rect 1489 532 1582 537
rect 345 522 462 527
rect 601 522 662 527
rect 713 522 830 527
rect 1145 522 1198 527
rect 1313 522 1342 527
rect 1337 517 1342 522
rect 1441 522 1470 527
rect 1633 522 1678 527
rect 1873 522 1982 527
rect 2081 522 2220 527
rect 1441 517 1446 522
rect 169 512 262 517
rect 609 512 638 517
rect 633 507 638 512
rect 737 512 766 517
rect 1337 512 1446 517
rect 1489 512 1598 517
rect 1649 512 1686 517
rect 1849 512 2030 517
rect 2081 512 2086 522
rect 737 507 742 512
rect 105 502 198 507
rect 225 502 270 507
rect 361 502 414 507
rect 633 502 742 507
rect 1609 502 1670 507
rect 1713 502 1822 507
rect 1945 502 1974 507
rect 2065 502 2102 507
rect 2113 502 2220 507
rect 2113 497 2118 502
rect 241 492 270 497
rect 409 492 566 497
rect 1777 492 1806 497
rect 1801 477 1806 492
rect 1977 492 2118 497
rect 1977 477 1982 492
rect 2001 482 2094 487
rect 1801 472 1982 477
rect 2017 472 2220 477
rect 257 432 390 437
rect 1473 432 1518 437
rect 321 422 366 427
rect 529 422 726 427
rect 153 412 238 417
rect 377 412 406 417
rect 529 407 534 422
rect 401 402 534 407
rect 721 407 726 422
rect 1769 422 1918 427
rect 1953 422 2006 427
rect 785 412 878 417
rect 937 412 1022 417
rect 1041 412 1142 417
rect 1321 412 1414 417
rect 1433 412 1558 417
rect 1577 412 1670 417
rect 1697 412 1726 417
rect 937 407 942 412
rect 721 402 742 407
rect 737 397 742 402
rect 817 402 942 407
rect 1017 407 1022 412
rect 1321 407 1326 412
rect 1017 402 1110 407
rect 1161 402 1278 407
rect 1297 402 1326 407
rect 1409 407 1414 412
rect 1577 407 1582 412
rect 1409 402 1582 407
rect 1665 407 1670 412
rect 1769 407 1774 422
rect 1665 402 1694 407
rect 1737 402 1774 407
rect 1913 407 1918 422
rect 1913 402 2094 407
rect 817 397 822 402
rect 1161 397 1166 402
rect 137 392 190 397
rect 369 392 398 397
rect 529 392 710 397
rect 737 392 822 397
rect 1065 392 1166 397
rect 1273 397 1278 402
rect 1273 392 1366 397
rect 1505 392 1686 397
rect 1785 392 1902 397
rect 673 382 678 392
rect 945 382 1046 387
rect 1353 382 1494 387
rect 1697 382 1758 387
rect 1833 382 2086 387
rect 1489 377 1702 382
rect 1177 372 1310 377
rect 1329 367 1446 372
rect 209 362 414 367
rect 561 362 606 367
rect 1033 362 1334 367
rect 1441 362 1686 367
rect 2073 362 2220 367
rect 409 352 614 357
rect 1113 352 1190 357
rect 1345 352 1430 357
rect 1921 352 1998 357
rect 2089 352 2118 357
rect 1185 347 1350 352
rect 145 342 246 347
rect 817 342 878 347
rect 1025 342 1070 347
rect 1137 342 1166 347
rect 1161 337 1166 342
rect 1369 342 1438 347
rect 1561 342 1590 347
rect 1769 342 1982 347
rect 2041 342 2110 347
rect 1369 337 1374 342
rect 1161 332 1374 337
rect 489 322 638 327
rect 1969 322 1998 327
rect 113 312 174 317
rect 257 312 446 317
rect 1025 312 1494 317
rect 1969 312 1974 322
rect 1993 317 1998 322
rect 2105 322 2220 327
rect 2105 317 2110 322
rect 1993 312 2110 317
rect 153 302 254 307
rect 377 302 406 307
rect 2129 302 2220 307
rect 1073 282 1206 287
rect 921 272 1030 277
rect 921 267 926 272
rect 137 262 190 267
rect 561 262 678 267
rect 897 262 926 267
rect 1025 267 1030 272
rect 1073 267 1078 282
rect 1025 262 1078 267
rect 1201 267 1206 282
rect 1249 272 1598 277
rect 1201 262 1230 267
rect 561 257 566 262
rect 537 252 566 257
rect 673 257 678 262
rect 1249 257 1254 272
rect 673 252 1254 257
rect 1593 257 1598 272
rect 1593 252 1622 257
rect 497 242 542 247
rect 553 242 662 247
rect 841 242 942 247
rect 1265 242 1510 247
rect 937 237 1054 242
rect 1153 237 1270 242
rect 73 232 118 237
rect 361 232 414 237
rect 1049 232 1158 237
rect 1353 227 1462 232
rect 1505 227 1510 242
rect 1633 242 1670 247
rect 1825 242 1894 247
rect 1633 227 1638 242
rect 1825 237 1830 242
rect 1801 232 1830 237
rect 1889 237 1894 242
rect 1889 232 2102 237
rect 97 222 134 227
rect 209 222 270 227
rect 425 222 1030 227
rect 1177 222 1222 227
rect 1273 222 1358 227
rect 1457 222 1486 227
rect 1505 222 1638 227
rect 1393 212 1478 217
rect 1841 212 1878 217
rect 705 202 822 207
rect 1713 202 1822 207
rect 705 197 710 202
rect 321 192 366 197
rect 401 192 710 197
rect 817 197 822 202
rect 817 192 846 197
rect 1761 192 1854 197
rect 1905 192 1958 197
rect 153 182 190 187
rect 721 182 814 187
rect 1081 182 1238 187
rect 1809 182 1974 187
rect 265 172 566 177
rect 721 172 750 177
rect 1249 172 1342 177
rect 785 167 878 172
rect 761 162 790 167
rect 873 162 902 167
rect 1001 162 1126 167
rect 2081 162 2220 167
rect 121 152 166 157
rect 201 152 278 157
rect 345 152 382 157
rect 569 152 806 157
rect 825 152 886 157
rect 1049 152 1262 157
rect 1473 152 1598 157
rect 121 142 286 147
rect 329 142 454 147
rect 465 142 566 147
rect 449 137 454 142
rect 561 137 566 142
rect 649 142 678 147
rect 785 142 822 147
rect 881 142 1046 147
rect 649 137 654 142
rect 1089 137 1094 147
rect 1857 142 2046 147
rect 449 132 542 137
rect 561 132 654 137
rect 985 132 1094 137
rect 761 127 934 132
rect 737 122 766 127
rect 929 122 958 127
rect 1417 122 1486 127
rect 249 112 358 117
rect 377 112 414 117
rect 505 112 582 117
rect 721 112 758 117
rect 793 112 838 117
rect 857 112 894 117
rect 1353 112 1438 117
rect 1545 112 1614 117
rect 273 102 302 107
rect 297 97 302 102
rect 377 102 406 107
rect 697 102 790 107
rect 1225 102 1374 107
rect 1409 102 1438 107
rect 377 97 382 102
rect 1433 97 1438 102
rect 1529 102 1558 107
rect 1529 97 1534 102
rect 297 92 382 97
rect 729 92 790 97
rect 1433 92 1534 97
rect 1777 82 1806 87
rect 1849 82 1878 87
rect 1905 82 1934 87
use top_module_VIA1  top_module_VIA1_0
timestamp 1681685098
transform 1 0 24 0 1 2017
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_1
timestamp 1681685098
transform 1 0 2194 0 1 2017
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_2
timestamp 1681685098
transform 1 0 48 0 1 1993
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_3
timestamp 1681685098
transform 1 0 2170 0 1 1993
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_0
timestamp 1681685098
transform 1 0 48 0 1 1970
box -10 -3 10 3
use M3_M2  M3_M2_13
timestamp 1681685098
transform 1 0 116 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_7
timestamp 1681685098
transform 1 0 196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1681685098
transform 1 0 116 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1681685098
transform 1 0 164 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_39
timestamp 1681685098
transform 1 0 196 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1681685098
transform 1 0 228 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_0
timestamp 1681685098
transform 1 0 236 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1681685098
transform 1 0 212 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1681685098
transform 1 0 244 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_15
timestamp 1681685098
transform 1 0 268 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_8
timestamp 1681685098
transform 1 0 268 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_16
timestamp 1681685098
transform 1 0 324 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_9
timestamp 1681685098
transform 1 0 324 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1681685098
transform 1 0 292 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_40
timestamp 1681685098
transform 1 0 324 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1681685098
transform 1 0 364 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_10
timestamp 1681685098
transform 1 0 436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1681685098
transform 1 0 356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1681685098
transform 1 0 396 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_41
timestamp 1681685098
transform 1 0 436 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_51
timestamp 1681685098
transform 1 0 452 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_42
timestamp 1681685098
transform 1 0 476 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1681685098
transform 1 0 516 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_1
timestamp 1681685098
transform 1 0 516 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_18
timestamp 1681685098
transform 1 0 540 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1681685098
transform 1 0 540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1681685098
transform 1 0 540 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_3
timestamp 1681685098
transform 1 0 572 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_12
timestamp 1681685098
transform 1 0 572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1681685098
transform 1 0 556 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_6
timestamp 1681685098
transform 1 0 628 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1681685098
transform 1 0 620 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_13
timestamp 1681685098
transform 1 0 620 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1681685098
transform 1 0 700 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1681685098
transform 1 0 716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1681685098
transform 1 0 708 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_7
timestamp 1681685098
transform 1 0 732 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1681685098
transform 1 0 780 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1681685098
transform 1 0 820 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_15
timestamp 1681685098
transform 1 0 804 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1681685098
transform 1 0 820 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1681685098
transform 1 0 780 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_43
timestamp 1681685098
transform 1 0 804 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_76
timestamp 1681685098
transform 1 0 820 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1681685098
transform 1 0 844 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1681685098
transform 1 0 876 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1681685098
transform 1 0 980 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1681685098
transform 1 0 956 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1681685098
transform 1 0 1004 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_19
timestamp 1681685098
transform 1 0 916 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1681685098
transform 1 0 916 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_20
timestamp 1681685098
transform 1 0 1012 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1681685098
transform 1 0 940 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1681685098
transform 1 0 996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1681685098
transform 1 0 1004 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1681685098
transform 1 0 1020 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1
timestamp 1681685098
transform 1 0 1068 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1681685098
transform 1 0 1052 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1681685098
transform 1 0 1044 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_45
timestamp 1681685098
transform 1 0 1044 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_3
timestamp 1681685098
transform 1 0 1100 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1681685098
transform 1 0 1092 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_9
timestamp 1681685098
transform 1 0 1116 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1681685098
transform 1 0 1108 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1681685098
transform 1 0 1100 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1681685098
transform 1 0 1156 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1681685098
transform 1 0 1140 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1681685098
transform 1 0 1220 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_23
timestamp 1681685098
transform 1 0 1188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1681685098
transform 1 0 1212 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_47
timestamp 1681685098
transform 1 0 1132 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_59
timestamp 1681685098
transform 1 0 1140 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_48
timestamp 1681685098
transform 1 0 1156 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_60
timestamp 1681685098
transform 1 0 1172 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_53
timestamp 1681685098
transform 1 0 1140 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1681685098
transform 1 0 1188 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1681685098
transform 1 0 1204 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1681685098
transform 1 0 1260 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1681685098
transform 1 0 1236 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1681685098
transform 1 0 1276 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_4
timestamp 1681685098
transform 1 0 1340 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1681685098
transform 1 0 1236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1681685098
transform 1 0 1252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1681685098
transform 1 0 1340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1681685098
transform 1 0 1276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1681685098
transform 1 0 1332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1681685098
transform 1 0 1236 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_54
timestamp 1681685098
transform 1 0 1340 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1681685098
transform 1 0 1332 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1681685098
transform 1 0 1380 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_28
timestamp 1681685098
transform 1 0 1380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1681685098
transform 1 0 1412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1681685098
transform 1 0 1436 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1681685098
transform 1 0 1436 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_78
timestamp 1681685098
transform 1 0 1436 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1681685098
transform 1 0 1452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1681685098
transform 1 0 1508 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_27
timestamp 1681685098
transform 1 0 1516 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_31
timestamp 1681685098
transform 1 0 1484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1681685098
transform 1 0 1492 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_50
timestamp 1681685098
transform 1 0 1492 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_33
timestamp 1681685098
transform 1 0 1516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1681685098
transform 1 0 1500 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_55
timestamp 1681685098
transform 1 0 1500 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1681685098
transform 1 0 1484 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1681685098
transform 1 0 1556 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_65
timestamp 1681685098
transform 1 0 1556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1681685098
transform 1 0 1548 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1681685098
transform 1 0 1580 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_51
timestamp 1681685098
transform 1 0 1588 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_80
timestamp 1681685098
transform 1 0 1580 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1681685098
transform 1 0 1572 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_56
timestamp 1681685098
transform 1 0 1580 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1681685098
transform 1 0 1668 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1681685098
transform 1 0 1660 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_6
timestamp 1681685098
transform 1 0 1668 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1681685098
transform 1 0 1660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1681685098
transform 1 0 1644 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_52
timestamp 1681685098
transform 1 0 1676 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1681685098
transform 1 0 1724 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1681685098
transform 1 0 1812 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_35
timestamp 1681685098
transform 1 0 1724 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1681685098
transform 1 0 1812 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1681685098
transform 1 0 1724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1681685098
transform 1 0 1732 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1681685098
transform 1 0 1764 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_61
timestamp 1681685098
transform 1 0 1716 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_37
timestamp 1681685098
transform 1 0 1828 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_62
timestamp 1681685098
transform 1 0 1828 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1681685098
transform 1 0 1852 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_38
timestamp 1681685098
transform 1 0 1860 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_37
timestamp 1681685098
transform 1 0 1868 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_39
timestamp 1681685098
transform 1 0 1884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1681685098
transform 1 0 1868 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1681685098
transform 1 0 1884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1681685098
transform 1 0 1884 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_63
timestamp 1681685098
transform 1 0 1884 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_40
timestamp 1681685098
transform 1 0 1916 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_32
timestamp 1681685098
transform 1 0 1932 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1681685098
transform 1 0 1980 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_41
timestamp 1681685098
transform 1 0 1932 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_38
timestamp 1681685098
transform 1 0 2028 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_42
timestamp 1681685098
transform 1 0 2036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1681685098
transform 1 0 1980 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1681685098
transform 1 0 2012 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_64
timestamp 1681685098
transform 1 0 1940 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1681685098
transform 1 0 1988 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1681685098
transform 1 0 2012 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1681685098
transform 1 0 2060 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_43
timestamp 1681685098
transform 1 0 2060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1681685098
transform 1 0 2068 0 1 1915
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_1
timestamp 1681685098
transform 1 0 2170 0 1 1970
box -10 -3 10 3
use top_module_VIA0  top_module_VIA0_2
timestamp 1681685098
transform 1 0 24 0 1 1870
box -10 -3 10 3
use FILL  FILL_0
timestamp 1681685098
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1
timestamp 1681685098
transform 1 0 80 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2
timestamp 1681685098
transform 1 0 88 0 -1 1970
box -8 -3 16 105
use FILL  FILL_3
timestamp 1681685098
transform 1 0 96 0 -1 1970
box -8 -3 16 105
use FILL  FILL_4
timestamp 1681685098
transform 1 0 104 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1681685098
transform -1 0 208 0 -1 1970
box -8 -3 104 105
use OR2X1  OR2X1_0
timestamp 1681685098
transform -1 0 240 0 -1 1970
box -8 -3 40 105
use FILL  FILL_5
timestamp 1681685098
transform 1 0 240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6
timestamp 1681685098
transform 1 0 248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7
timestamp 1681685098
transform 1 0 256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_8
timestamp 1681685098
transform 1 0 264 0 -1 1970
box -8 -3 16 105
use XNOR2X1  XNOR2X1_0
timestamp 1681685098
transform -1 0 328 0 -1 1970
box -8 -3 64 105
use FILL  FILL_9
timestamp 1681685098
transform 1 0 328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_10
timestamp 1681685098
transform 1 0 336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_11
timestamp 1681685098
transform 1 0 344 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1681685098
transform -1 0 448 0 -1 1970
box -8 -3 104 105
use FILL  FILL_12
timestamp 1681685098
transform 1 0 448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_13
timestamp 1681685098
transform 1 0 456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_14
timestamp 1681685098
transform 1 0 464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_15
timestamp 1681685098
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use OR2X1  OR2X1_1
timestamp 1681685098
transform -1 0 512 0 -1 1970
box -8 -3 40 105
use FILL  FILL_16
timestamp 1681685098
transform 1 0 512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_17
timestamp 1681685098
transform 1 0 520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_18
timestamp 1681685098
transform 1 0 528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_19
timestamp 1681685098
transform 1 0 536 0 -1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1681685098
transform -1 0 568 0 -1 1970
box -8 -3 32 105
use XNOR2X1  XNOR2X1_1
timestamp 1681685098
transform -1 0 624 0 -1 1970
box -8 -3 64 105
use FILL  FILL_20
timestamp 1681685098
transform 1 0 624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_21
timestamp 1681685098
transform 1 0 632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_22
timestamp 1681685098
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_23
timestamp 1681685098
transform 1 0 648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_24
timestamp 1681685098
transform 1 0 656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_25
timestamp 1681685098
transform 1 0 664 0 -1 1970
box -8 -3 16 105
use OR2X1  OR2X1_2
timestamp 1681685098
transform -1 0 704 0 -1 1970
box -8 -3 40 105
use FILL  FILL_26
timestamp 1681685098
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_27
timestamp 1681685098
transform 1 0 712 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1681685098
transform -1 0 816 0 -1 1970
box -8 -3 104 105
use OAI21X1  OAI21X1_0
timestamp 1681685098
transform -1 0 848 0 -1 1970
box -8 -3 34 105
use FILL  FILL_28
timestamp 1681685098
transform 1 0 848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_29
timestamp 1681685098
transform 1 0 856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_30
timestamp 1681685098
transform 1 0 864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_31
timestamp 1681685098
transform 1 0 872 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1681685098
transform 1 0 880 0 -1 1970
box -9 -3 26 105
use FILL  FILL_32
timestamp 1681685098
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1681685098
transform 1 0 904 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_1
timestamp 1681685098
transform -1 0 1016 0 -1 1970
box -9 -3 26 105
use FILL  FILL_33
timestamp 1681685098
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_34
timestamp 1681685098
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_35
timestamp 1681685098
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use XNOR2X1  XNOR2X1_2
timestamp 1681685098
transform -1 0 1096 0 -1 1970
box -8 -3 64 105
use FILL  FILL_36
timestamp 1681685098
transform 1 0 1096 0 -1 1970
box -8 -3 16 105
use OR2X1  OR2X1_3
timestamp 1681685098
transform 1 0 1104 0 -1 1970
box -8 -3 40 105
use XNOR2X1  XNOR2X1_3
timestamp 1681685098
transform 1 0 1136 0 -1 1970
box -8 -3 64 105
use INVX2  INVX2_2
timestamp 1681685098
transform 1 0 1192 0 -1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_1
timestamp 1681685098
transform 1 0 1208 0 -1 1970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1681685098
transform 1 0 1240 0 -1 1970
box -8 -3 104 105
use OR2X1  OR2X1_4
timestamp 1681685098
transform 1 0 1336 0 -1 1970
box -8 -3 40 105
use FILL  FILL_37
timestamp 1681685098
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use XNOR2X1  XNOR2X1_4
timestamp 1681685098
transform 1 0 1376 0 -1 1970
box -8 -3 64 105
use FILL  FILL_38
timestamp 1681685098
transform 1 0 1432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_39
timestamp 1681685098
transform 1 0 1440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_40
timestamp 1681685098
transform 1 0 1448 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1681685098
transform -1 0 1488 0 -1 1970
box -8 -3 34 105
use INVX2  INVX2_3
timestamp 1681685098
transform 1 0 1488 0 -1 1970
box -9 -3 26 105
use OR2X1  OR2X1_5
timestamp 1681685098
transform 1 0 1504 0 -1 1970
box -8 -3 40 105
use FILL  FILL_41
timestamp 1681685098
transform 1 0 1536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_42
timestamp 1681685098
transform 1 0 1544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_43
timestamp 1681685098
transform 1 0 1552 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1681685098
transform -1 0 1592 0 -1 1970
box -8 -3 40 105
use FILL  FILL_44
timestamp 1681685098
transform 1 0 1592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_45
timestamp 1681685098
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_46
timestamp 1681685098
transform 1 0 1608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_47
timestamp 1681685098
transform 1 0 1616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_48
timestamp 1681685098
transform 1 0 1624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_49
timestamp 1681685098
transform 1 0 1632 0 -1 1970
box -8 -3 16 105
use OR2X1  OR2X1_6
timestamp 1681685098
transform -1 0 1672 0 -1 1970
box -8 -3 40 105
use M3_M2  M3_M2_67
timestamp 1681685098
transform 1 0 1724 0 1 1875
box -3 -3 3 3
use XNOR2X1  XNOR2X1_5
timestamp 1681685098
transform 1 0 1672 0 -1 1970
box -8 -3 64 105
use M3_M2  M3_M2_68
timestamp 1681685098
transform 1 0 1764 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_5
timestamp 1681685098
transform -1 0 1824 0 -1 1970
box -8 -3 104 105
use FILL  FILL_50
timestamp 1681685098
transform 1 0 1824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_51
timestamp 1681685098
transform 1 0 1832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_52
timestamp 1681685098
transform 1 0 1840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_53
timestamp 1681685098
transform 1 0 1848 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1681685098
transform 1 0 1856 0 -1 1970
box -8 -3 34 105
use INVX2  INVX2_4
timestamp 1681685098
transform -1 0 1904 0 -1 1970
box -9 -3 26 105
use FILL  FILL_54
timestamp 1681685098
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_55
timestamp 1681685098
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1681685098
transform 1 0 1920 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_5
timestamp 1681685098
transform 1 0 2016 0 -1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_4
timestamp 1681685098
transform 1 0 2032 0 -1 1970
box -8 -3 34 105
use FILL  FILL_56
timestamp 1681685098
transform 1 0 2064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_57
timestamp 1681685098
transform 1 0 2072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_58
timestamp 1681685098
transform 1 0 2080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_59
timestamp 1681685098
transform 1 0 2088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_60
timestamp 1681685098
transform 1 0 2096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_61
timestamp 1681685098
transform 1 0 2104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_62
timestamp 1681685098
transform 1 0 2112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_63
timestamp 1681685098
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_64
timestamp 1681685098
transform 1 0 2128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_65
timestamp 1681685098
transform 1 0 2136 0 -1 1970
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_3
timestamp 1681685098
transform 1 0 2194 0 1 1870
box -10 -3 10 3
use M3_M2  M3_M2_120
timestamp 1681685098
transform 1 0 84 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_94
timestamp 1681685098
transform 1 0 100 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1681685098
transform 1 0 124 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1681685098
transform 1 0 164 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1681685098
transform 1 0 172 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1681685098
transform 1 0 180 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_95
timestamp 1681685098
transform 1 0 196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1681685098
transform 1 0 220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1681685098
transform 1 0 196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1681685098
transform 1 0 204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1681685098
transform 1 0 212 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_103
timestamp 1681685098
transform 1 0 196 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1681685098
transform 1 0 196 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_166
timestamp 1681685098
transform 1 0 220 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_122
timestamp 1681685098
transform 1 0 220 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_130
timestamp 1681685098
transform 1 0 244 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_123
timestamp 1681685098
transform 1 0 268 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1681685098
transform 1 0 300 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_97
timestamp 1681685098
transform 1 0 300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1681685098
transform 1 0 284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1681685098
transform 1 0 292 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_104
timestamp 1681685098
transform 1 0 300 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_85
timestamp 1681685098
transform 1 0 332 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_79
timestamp 1681685098
transform 1 0 372 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_98
timestamp 1681685098
transform 1 0 348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1681685098
transform 1 0 364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1681685098
transform 1 0 356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1681685098
transform 1 0 380 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_105
timestamp 1681685098
transform 1 0 364 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1681685098
transform 1 0 380 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1681685098
transform 1 0 412 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_100
timestamp 1681685098
transform 1 0 412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1681685098
transform 1 0 388 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_124
timestamp 1681685098
transform 1 0 356 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1681685098
transform 1 0 388 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_135
timestamp 1681685098
transform 1 0 444 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_107
timestamp 1681685098
transform 1 0 444 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_86
timestamp 1681685098
transform 1 0 564 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1681685098
transform 1 0 524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1681685098
transform 1 0 564 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_87
timestamp 1681685098
transform 1 0 572 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_136
timestamp 1681685098
transform 1 0 476 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1681685098
transform 1 0 564 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_108
timestamp 1681685098
transform 1 0 524 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1681685098
transform 1 0 564 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_138
timestamp 1681685098
transform 1 0 588 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_110
timestamp 1681685098
transform 1 0 636 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1681685098
transform 1 0 652 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_139
timestamp 1681685098
transform 1 0 652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1681685098
transform 1 0 668 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_111
timestamp 1681685098
transform 1 0 668 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_141
timestamp 1681685098
transform 1 0 684 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1681685098
transform 1 0 700 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_97
timestamp 1681685098
transform 1 0 700 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_104
timestamp 1681685098
transform 1 0 772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1681685098
transform 1 0 780 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_98
timestamp 1681685098
transform 1 0 788 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1681685098
transform 1 0 780 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_105
timestamp 1681685098
transform 1 0 820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1681685098
transform 1 0 844 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_73
timestamp 1681685098
transform 1 0 884 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_106
timestamp 1681685098
transform 1 0 884 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_99
timestamp 1681685098
transform 1 0 876 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_143
timestamp 1681685098
transform 1 0 900 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_69
timestamp 1681685098
transform 1 0 924 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1681685098
transform 1 0 916 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_87
timestamp 1681685098
transform 1 0 916 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_113
timestamp 1681685098
transform 1 0 892 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1681685098
transform 1 0 908 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_107
timestamp 1681685098
transform 1 0 924 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1681685098
transform 1 0 932 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_100
timestamp 1681685098
transform 1 0 940 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1681685098
transform 1 0 964 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_108
timestamp 1681685098
transform 1 0 964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1681685098
transform 1 0 956 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_126
timestamp 1681685098
transform 1 0 956 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1681685098
transform 1 0 1020 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1681685098
transform 1 0 1004 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1681685098
transform 1 0 980 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_109
timestamp 1681685098
transform 1 0 1012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1681685098
transform 1 0 1060 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1681685098
transform 1 0 980 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_115
timestamp 1681685098
transform 1 0 980 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_111
timestamp 1681685098
transform 1 0 1092 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1681685098
transform 1 0 1076 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1681685098
transform 1 0 1068 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_75
timestamp 1681685098
transform 1 0 1156 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_88
timestamp 1681685098
transform 1 0 1148 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_90
timestamp 1681685098
transform 1 0 1148 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1681685098
transform 1 0 1140 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1681685098
transform 1 0 1156 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1681685098
transform 1 0 1180 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_112
timestamp 1681685098
transform 1 0 1180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1681685098
transform 1 0 1172 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_76
timestamp 1681685098
transform 1 0 1204 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_113
timestamp 1681685098
transform 1 0 1196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1681685098
transform 1 0 1212 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_128
timestamp 1681685098
transform 1 0 1212 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1681685098
transform 1 0 1252 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1681685098
transform 1 0 1284 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1681685098
transform 1 0 1236 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1681685098
transform 1 0 1228 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_114
timestamp 1681685098
transform 1 0 1252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1681685098
transform 1 0 1260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1681685098
transform 1 0 1316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1681685098
transform 1 0 1236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1681685098
transform 1 0 1228 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_117
timestamp 1681685098
transform 1 0 1244 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_151
timestamp 1681685098
transform 1 0 1340 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_118
timestamp 1681685098
transform 1 0 1340 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1681685098
transform 1 0 1260 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_89
timestamp 1681685098
transform 1 0 1372 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_91
timestamp 1681685098
transform 1 0 1372 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_90
timestamp 1681685098
transform 1 0 1396 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1681685098
transform 1 0 1412 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_119
timestamp 1681685098
transform 1 0 1420 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_117
timestamp 1681685098
transform 1 0 1436 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_102
timestamp 1681685098
transform 1 0 1548 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_153
timestamp 1681685098
transform 1 0 1572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1681685098
transform 1 0 1564 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_130
timestamp 1681685098
transform 1 0 1564 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_172
timestamp 1681685098
transform 1 0 1588 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_131
timestamp 1681685098
transform 1 0 1612 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_118
timestamp 1681685098
transform 1 0 1668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1681685098
transform 1 0 1676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1681685098
transform 1 0 1644 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1681685098
transform 1 0 1652 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_92
timestamp 1681685098
transform 1 0 1684 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_156
timestamp 1681685098
transform 1 0 1684 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1681685098
transform 1 0 1716 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_93
timestamp 1681685098
transform 1 0 1732 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_158
timestamp 1681685098
transform 1 0 1732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1681685098
transform 1 0 1780 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_94
timestamp 1681685098
transform 1 0 1780 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_159
timestamp 1681685098
transform 1 0 1756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1681685098
transform 1 0 1764 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1681685098
transform 1 0 1948 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1681685098
transform 1 0 1884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1681685098
transform 1 0 1932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1681685098
transform 1 0 1940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1681685098
transform 1 0 1852 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_95
timestamp 1681685098
transform 1 0 1948 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_162
timestamp 1681685098
transform 1 0 1980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1681685098
transform 1 0 1988 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_85
timestamp 1681685098
transform 1 0 2036 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_93
timestamp 1681685098
transform 1 0 2044 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1681685098
transform 1 0 2036 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_96
timestamp 1681685098
transform 1 0 2044 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_164
timestamp 1681685098
transform 1 0 2044 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_86
timestamp 1681685098
transform 1 0 2060 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_124
timestamp 1681685098
transform 1 0 2068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1681685098
transform 1 0 2060 0 1 1805
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_4
timestamp 1681685098
transform 1 0 48 0 1 1770
box -10 -3 10 3
use FILL  FILL_66
timestamp 1681685098
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_68
timestamp 1681685098
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_70
timestamp 1681685098
transform 1 0 88 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_6
timestamp 1681685098
transform -1 0 112 0 1 1770
box -9 -3 26 105
use FILL  FILL_71
timestamp 1681685098
transform 1 0 112 0 1 1770
box -8 -3 16 105
use FILL  FILL_72
timestamp 1681685098
transform 1 0 120 0 1 1770
box -8 -3 16 105
use FILL  FILL_74
timestamp 1681685098
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_76
timestamp 1681685098
transform 1 0 136 0 1 1770
box -8 -3 16 105
use FILL  FILL_78
timestamp 1681685098
transform 1 0 144 0 1 1770
box -8 -3 16 105
use FILL  FILL_80
timestamp 1681685098
transform 1 0 152 0 1 1770
box -8 -3 16 105
use FILL  FILL_82
timestamp 1681685098
transform 1 0 160 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1681685098
transform -1 0 200 0 1 1770
box -8 -3 34 105
use NOR2X1  NOR2X1_0
timestamp 1681685098
transform -1 0 224 0 1 1770
box -8 -3 32 105
use INVX2  INVX2_7
timestamp 1681685098
transform -1 0 240 0 1 1770
box -9 -3 26 105
use FILL  FILL_83
timestamp 1681685098
transform 1 0 240 0 1 1770
box -8 -3 16 105
use FILL  FILL_84
timestamp 1681685098
transform 1 0 248 0 1 1770
box -8 -3 16 105
use FILL  FILL_85
timestamp 1681685098
transform 1 0 256 0 1 1770
box -8 -3 16 105
use FILL  FILL_86
timestamp 1681685098
transform 1 0 264 0 1 1770
box -8 -3 16 105
use FILL  FILL_87
timestamp 1681685098
transform 1 0 272 0 1 1770
box -8 -3 16 105
use FILL  FILL_88
timestamp 1681685098
transform 1 0 280 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1681685098
transform 1 0 288 0 1 1770
box -8 -3 32 105
use FILL  FILL_89
timestamp 1681685098
transform 1 0 312 0 1 1770
box -8 -3 16 105
use FILL  FILL_95
timestamp 1681685098
transform 1 0 320 0 1 1770
box -8 -3 16 105
use FILL  FILL_97
timestamp 1681685098
transform 1 0 328 0 1 1770
box -8 -3 16 105
use FILL  FILL_99
timestamp 1681685098
transform 1 0 336 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_8
timestamp 1681685098
transform -1 0 360 0 1 1770
box -9 -3 26 105
use OR2X1  OR2X1_8
timestamp 1681685098
transform -1 0 392 0 1 1770
box -8 -3 40 105
use XNOR2X1  XNOR2X1_7
timestamp 1681685098
transform -1 0 448 0 1 1770
box -8 -3 64 105
use FILL  FILL_100
timestamp 1681685098
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_101
timestamp 1681685098
transform 1 0 456 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1681685098
transform 1 0 464 0 1 1770
box -8 -3 104 105
use OAI21X1  OAI21X1_7
timestamp 1681685098
transform -1 0 592 0 1 1770
box -8 -3 34 105
use FILL  FILL_102
timestamp 1681685098
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_122
timestamp 1681685098
transform 1 0 600 0 1 1770
box -8 -3 16 105
use FILL  FILL_124
timestamp 1681685098
transform 1 0 608 0 1 1770
box -8 -3 16 105
use FILL  FILL_126
timestamp 1681685098
transform 1 0 616 0 1 1770
box -8 -3 16 105
use FILL  FILL_127
timestamp 1681685098
transform 1 0 624 0 1 1770
box -8 -3 16 105
use FILL  FILL_128
timestamp 1681685098
transform 1 0 632 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_10
timestamp 1681685098
transform -1 0 656 0 1 1770
box -9 -3 26 105
use NOR2X1  NOR2X1_1
timestamp 1681685098
transform 1 0 656 0 1 1770
box -8 -3 32 105
use FILL  FILL_129
timestamp 1681685098
transform 1 0 680 0 1 1770
box -8 -3 16 105
use FILL  FILL_133
timestamp 1681685098
transform 1 0 688 0 1 1770
box -8 -3 16 105
use FILL  FILL_135
timestamp 1681685098
transform 1 0 696 0 1 1770
box -8 -3 16 105
use FILL  FILL_137
timestamp 1681685098
transform 1 0 704 0 1 1770
box -8 -3 16 105
use FILL  FILL_138
timestamp 1681685098
transform 1 0 712 0 1 1770
box -8 -3 16 105
use FILL  FILL_139
timestamp 1681685098
transform 1 0 720 0 1 1770
box -8 -3 16 105
use FILL  FILL_140
timestamp 1681685098
transform 1 0 728 0 1 1770
box -8 -3 16 105
use FILL  FILL_141
timestamp 1681685098
transform 1 0 736 0 1 1770
box -8 -3 16 105
use FILL  FILL_142
timestamp 1681685098
transform 1 0 744 0 1 1770
box -8 -3 16 105
use FILL  FILL_143
timestamp 1681685098
transform 1 0 752 0 1 1770
box -8 -3 16 105
use FILL  FILL_144
timestamp 1681685098
transform 1 0 760 0 1 1770
box -8 -3 16 105
use AOI21X1  AOI21X1_0
timestamp 1681685098
transform 1 0 768 0 1 1770
box -7 -3 39 105
use FILL  FILL_145
timestamp 1681685098
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_146
timestamp 1681685098
transform 1 0 808 0 1 1770
box -8 -3 16 105
use FILL  FILL_147
timestamp 1681685098
transform 1 0 816 0 1 1770
box -8 -3 16 105
use FILL  FILL_148
timestamp 1681685098
transform 1 0 824 0 1 1770
box -8 -3 16 105
use FILL  FILL_150
timestamp 1681685098
transform 1 0 832 0 1 1770
box -8 -3 16 105
use FILL  FILL_151
timestamp 1681685098
transform 1 0 840 0 1 1770
box -8 -3 16 105
use FILL  FILL_152
timestamp 1681685098
transform 1 0 848 0 1 1770
box -8 -3 16 105
use FILL  FILL_153
timestamp 1681685098
transform 1 0 856 0 1 1770
box -8 -3 16 105
use FILL  FILL_156
timestamp 1681685098
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_158
timestamp 1681685098
transform 1 0 872 0 1 1770
box -8 -3 16 105
use AOI21X1  AOI21X1_1
timestamp 1681685098
transform -1 0 912 0 1 1770
box -7 -3 39 105
use FILL  FILL_159
timestamp 1681685098
transform 1 0 912 0 1 1770
box -8 -3 16 105
use FILL  FILL_160
timestamp 1681685098
transform 1 0 920 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_11
timestamp 1681685098
transform -1 0 960 0 1 1770
box -8 -3 34 105
use FILL  FILL_161
timestamp 1681685098
transform 1 0 960 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1681685098
transform 1 0 968 0 1 1770
box -8 -3 104 105
use OR2X1  OR2X1_11
timestamp 1681685098
transform 1 0 1064 0 1 1770
box -8 -3 40 105
use FILL  FILL_171
timestamp 1681685098
transform 1 0 1096 0 1 1770
box -8 -3 16 105
use FILL  FILL_183
timestamp 1681685098
transform 1 0 1104 0 1 1770
box -8 -3 16 105
use FILL  FILL_185
timestamp 1681685098
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_187
timestamp 1681685098
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use FILL  FILL_188
timestamp 1681685098
transform 1 0 1128 0 1 1770
box -8 -3 16 105
use FILL  FILL_189
timestamp 1681685098
transform 1 0 1136 0 1 1770
box -8 -3 16 105
use FILL  FILL_190
timestamp 1681685098
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_3
timestamp 1681685098
transform -1 0 1176 0 1 1770
box -8 -3 32 105
use FILL  FILL_191
timestamp 1681685098
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_197
timestamp 1681685098
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_199
timestamp 1681685098
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_14
timestamp 1681685098
transform -1 0 1216 0 1 1770
box -9 -3 26 105
use FILL  FILL_200
timestamp 1681685098
transform 1 0 1216 0 1 1770
box -8 -3 16 105
use OR2X1  OR2X1_12
timestamp 1681685098
transform 1 0 1224 0 1 1770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1681685098
transform -1 0 1352 0 1 1770
box -8 -3 104 105
use FILL  FILL_201
timestamp 1681685098
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use FILL  FILL_215
timestamp 1681685098
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use FILL  FILL_217
timestamp 1681685098
transform 1 0 1368 0 1 1770
box -8 -3 16 105
use FILL  FILL_219
timestamp 1681685098
transform 1 0 1376 0 1 1770
box -8 -3 16 105
use FILL  FILL_221
timestamp 1681685098
transform 1 0 1384 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1681685098
transform -1 0 1416 0 1 1770
box -8 -3 32 105
use FILL  FILL_222
timestamp 1681685098
transform 1 0 1416 0 1 1770
box -8 -3 16 105
use FILL  FILL_223
timestamp 1681685098
transform 1 0 1424 0 1 1770
box -8 -3 16 105
use FILL  FILL_224
timestamp 1681685098
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_225
timestamp 1681685098
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use FILL  FILL_226
timestamp 1681685098
transform 1 0 1448 0 1 1770
box -8 -3 16 105
use FILL  FILL_227
timestamp 1681685098
transform 1 0 1456 0 1 1770
box -8 -3 16 105
use FILL  FILL_228
timestamp 1681685098
transform 1 0 1464 0 1 1770
box -8 -3 16 105
use FILL  FILL_229
timestamp 1681685098
transform 1 0 1472 0 1 1770
box -8 -3 16 105
use FILL  FILL_230
timestamp 1681685098
transform 1 0 1480 0 1 1770
box -8 -3 16 105
use FILL  FILL_231
timestamp 1681685098
transform 1 0 1488 0 1 1770
box -8 -3 16 105
use FILL  FILL_232
timestamp 1681685098
transform 1 0 1496 0 1 1770
box -8 -3 16 105
use FILL  FILL_233
timestamp 1681685098
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_234
timestamp 1681685098
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_235
timestamp 1681685098
transform 1 0 1520 0 1 1770
box -8 -3 16 105
use FILL  FILL_236
timestamp 1681685098
transform 1 0 1528 0 1 1770
box -8 -3 16 105
use FILL  FILL_237
timestamp 1681685098
transform 1 0 1536 0 1 1770
box -8 -3 16 105
use FILL  FILL_238
timestamp 1681685098
transform 1 0 1544 0 1 1770
box -8 -3 16 105
use FILL  FILL_239
timestamp 1681685098
transform 1 0 1552 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_3
timestamp 1681685098
transform 1 0 1560 0 1 1770
box -8 -3 32 105
use FILL  FILL_240
timestamp 1681685098
transform 1 0 1584 0 1 1770
box -8 -3 16 105
use FILL  FILL_241
timestamp 1681685098
transform 1 0 1592 0 1 1770
box -8 -3 16 105
use FILL  FILL_242
timestamp 1681685098
transform 1 0 1600 0 1 1770
box -8 -3 16 105
use FILL  FILL_243
timestamp 1681685098
transform 1 0 1608 0 1 1770
box -8 -3 16 105
use FILL  FILL_244
timestamp 1681685098
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_245
timestamp 1681685098
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use FILL  FILL_246
timestamp 1681685098
transform 1 0 1632 0 1 1770
box -8 -3 16 105
use OR2X1  OR2X1_13
timestamp 1681685098
transform 1 0 1640 0 1 1770
box -8 -3 40 105
use FILL  FILL_247
timestamp 1681685098
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_15
timestamp 1681685098
transform 1 0 1680 0 1 1770
box -9 -3 26 105
use FILL  FILL_248
timestamp 1681685098
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use FILL  FILL_249
timestamp 1681685098
transform 1 0 1704 0 1 1770
box -8 -3 16 105
use FILL  FILL_250
timestamp 1681685098
transform 1 0 1712 0 1 1770
box -8 -3 16 105
use FILL  FILL_251
timestamp 1681685098
transform 1 0 1720 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_14
timestamp 1681685098
transform 1 0 1728 0 1 1770
box -8 -3 34 105
use NAND2X1  NAND2X1_5
timestamp 1681685098
transform 1 0 1760 0 1 1770
box -8 -3 32 105
use FILL  FILL_259
timestamp 1681685098
transform 1 0 1784 0 1 1770
box -8 -3 16 105
use FILL  FILL_261
timestamp 1681685098
transform 1 0 1792 0 1 1770
box -8 -3 16 105
use FILL  FILL_263
timestamp 1681685098
transform 1 0 1800 0 1 1770
box -8 -3 16 105
use FILL  FILL_265
timestamp 1681685098
transform 1 0 1808 0 1 1770
box -8 -3 16 105
use FILL  FILL_267
timestamp 1681685098
transform 1 0 1816 0 1 1770
box -8 -3 16 105
use FILL  FILL_269
timestamp 1681685098
transform 1 0 1824 0 1 1770
box -8 -3 16 105
use FILL  FILL_271
timestamp 1681685098
transform 1 0 1832 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1681685098
transform 1 0 1840 0 1 1770
box -8 -3 104 105
use FILL  FILL_273
timestamp 1681685098
transform 1 0 1936 0 1 1770
box -8 -3 16 105
use FILL  FILL_283
timestamp 1681685098
transform 1 0 1944 0 1 1770
box -8 -3 16 105
use FILL  FILL_284
timestamp 1681685098
transform 1 0 1952 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_7
timestamp 1681685098
transform -1 0 1984 0 1 1770
box -8 -3 32 105
use XNOR2X1  XNOR2X1_11
timestamp 1681685098
transform 1 0 1984 0 1 1770
box -8 -3 64 105
use NAND2X1  NAND2X1_8
timestamp 1681685098
transform -1 0 2064 0 1 1770
box -8 -3 32 105
use FILL  FILL_285
timestamp 1681685098
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_288
timestamp 1681685098
transform 1 0 2072 0 1 1770
box -8 -3 16 105
use FILL  FILL_290
timestamp 1681685098
transform 1 0 2080 0 1 1770
box -8 -3 16 105
use FILL  FILL_292
timestamp 1681685098
transform 1 0 2088 0 1 1770
box -8 -3 16 105
use FILL  FILL_294
timestamp 1681685098
transform 1 0 2096 0 1 1770
box -8 -3 16 105
use FILL  FILL_296
timestamp 1681685098
transform 1 0 2104 0 1 1770
box -8 -3 16 105
use FILL  FILL_298
timestamp 1681685098
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use FILL  FILL_300
timestamp 1681685098
transform 1 0 2120 0 1 1770
box -8 -3 16 105
use FILL  FILL_302
timestamp 1681685098
transform 1 0 2128 0 1 1770
box -8 -3 16 105
use FILL  FILL_304
timestamp 1681685098
transform 1 0 2136 0 1 1770
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_5
timestamp 1681685098
transform 1 0 2170 0 1 1770
box -10 -3 10 3
use M2_M1  M2_M1_180
timestamp 1681685098
transform 1 0 84 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1681685098
transform 1 0 116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1681685098
transform 1 0 100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1681685098
transform 1 0 124 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1681685098
transform 1 0 132 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1681685098
transform 1 0 156 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_132
timestamp 1681685098
transform 1 0 196 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_174
timestamp 1681685098
transform 1 0 188 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1681685098
transform 1 0 196 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_133
timestamp 1681685098
transform 1 0 228 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_183
timestamp 1681685098
transform 1 0 268 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1681685098
transform 1 0 284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1681685098
transform 1 0 236 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_163
timestamp 1681685098
transform 1 0 212 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1681685098
transform 1 0 276 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_243
timestamp 1681685098
transform 1 0 284 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1681685098
transform 1 0 276 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_171
timestamp 1681685098
transform 1 0 284 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1681685098
transform 1 0 324 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_244
timestamp 1681685098
transform 1 0 324 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1681685098
transform 1 0 348 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_172
timestamp 1681685098
transform 1 0 348 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1681685098
transform 1 0 364 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_185
timestamp 1681685098
transform 1 0 364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1681685098
transform 1 0 388 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1681685098
transform 1 0 396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1681685098
transform 1 0 428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1681685098
transform 1 0 436 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_173
timestamp 1681685098
transform 1 0 436 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1681685098
transform 1 0 460 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_175
timestamp 1681685098
transform 1 0 484 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1681685098
transform 1 0 460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1681685098
transform 1 0 476 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_148
timestamp 1681685098
transform 1 0 484 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1681685098
transform 1 0 484 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_190
timestamp 1681685098
transform 1 0 556 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_155
timestamp 1681685098
transform 1 0 556 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1681685098
transform 1 0 588 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1681685098
transform 1 0 580 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_247
timestamp 1681685098
transform 1 0 580 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1681685098
transform 1 0 620 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1681685098
transform 1 0 644 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1681685098
transform 1 0 660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1681685098
transform 1 0 652 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1681685098
transform 1 0 636 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_175
timestamp 1681685098
transform 1 0 652 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_176
timestamp 1681685098
transform 1 0 708 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1681685098
transform 1 0 716 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_157
timestamp 1681685098
transform 1 0 716 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1681685098
transform 1 0 772 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_192
timestamp 1681685098
transform 1 0 788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1681685098
transform 1 0 796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1681685098
transform 1 0 732 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_158
timestamp 1681685098
transform 1 0 756 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_224
timestamp 1681685098
transform 1 0 772 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_165
timestamp 1681685098
transform 1 0 772 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1681685098
transform 1 0 828 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_194
timestamp 1681685098
transform 1 0 820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1681685098
transform 1 0 812 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1681685098
transform 1 0 796 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_176
timestamp 1681685098
transform 1 0 812 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1681685098
transform 1 0 796 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_195
timestamp 1681685098
transform 1 0 852 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1681685098
transform 1 0 908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1681685098
transform 1 0 900 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_178
timestamp 1681685098
transform 1 0 900 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_250
timestamp 1681685098
transform 1 0 924 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_149
timestamp 1681685098
transform 1 0 964 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_251
timestamp 1681685098
transform 1 0 964 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1681685098
transform 1 0 1012 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1681685098
transform 1 0 1004 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_145
timestamp 1681685098
transform 1 0 1044 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_198
timestamp 1681685098
transform 1 0 1044 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1681685098
transform 1 0 1052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1681685098
transform 1 0 1124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1681685098
transform 1 0 1132 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_166
timestamp 1681685098
transform 1 0 1124 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1681685098
transform 1 0 1148 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_200
timestamp 1681685098
transform 1 0 1156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1681685098
transform 1 0 1156 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1681685098
transform 1 0 1180 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_151
timestamp 1681685098
transform 1 0 1196 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_229
timestamp 1681685098
transform 1 0 1204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1681685098
transform 1 0 1196 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_167
timestamp 1681685098
transform 1 0 1204 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1681685098
transform 1 0 1244 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_201
timestamp 1681685098
transform 1 0 1236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1681685098
transform 1 0 1244 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_152
timestamp 1681685098
transform 1 0 1284 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_203
timestamp 1681685098
transform 1 0 1292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1681685098
transform 1 0 1284 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1681685098
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_134
timestamp 1681685098
transform 1 0 1396 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_254
timestamp 1681685098
transform 1 0 1388 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_135
timestamp 1681685098
transform 1 0 1428 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_205
timestamp 1681685098
transform 1 0 1420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1681685098
transform 1 0 1516 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_137
timestamp 1681685098
transform 1 0 1652 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1681685098
transform 1 0 1676 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_207
timestamp 1681685098
transform 1 0 1612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1681685098
transform 1 0 1452 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1681685098
transform 1 0 1500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1681685098
transform 1 0 1556 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_159
timestamp 1681685098
transform 1 0 1588 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_234
timestamp 1681685098
transform 1 0 1596 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1681685098
transform 1 0 1604 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1681685098
transform 1 0 1668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1681685098
transform 1 0 1676 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1681685098
transform 1 0 1652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1681685098
transform 1 0 1724 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_153
timestamp 1681685098
transform 1 0 1732 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1681685098
transform 1 0 1724 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_237
timestamp 1681685098
transform 1 0 1772 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1681685098
transform 1 0 1780 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1681685098
transform 1 0 1796 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1681685098
transform 1 0 1852 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_154
timestamp 1681685098
transform 1 0 1892 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_212
timestamp 1681685098
transform 1 0 1900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1681685098
transform 1 0 1908 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1681685098
transform 1 0 1932 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_168
timestamp 1681685098
transform 1 0 1932 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1681685098
transform 1 0 1972 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1681685098
transform 1 0 1988 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_178
timestamp 1681685098
transform 1 0 1972 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1681685098
transform 1 0 1964 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1681685098
transform 1 0 1972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1681685098
transform 1 0 1980 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_169
timestamp 1681685098
transform 1 0 1972 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_179
timestamp 1681685098
transform 1 0 2036 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1681685098
transform 1 0 2044 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_161
timestamp 1681685098
transform 1 0 2044 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_241
timestamp 1681685098
transform 1 0 2060 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_170
timestamp 1681685098
transform 1 0 2036 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1681685098
transform 1 0 2124 0 1 1725
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_6
timestamp 1681685098
transform 1 0 24 0 1 1670
box -10 -3 10 3
use FILL  FILL_67
timestamp 1681685098
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_69
timestamp 1681685098
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1681685098
transform 1 0 88 0 -1 1770
box -8 -3 34 105
use FILL  FILL_73
timestamp 1681685098
transform 1 0 120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_75
timestamp 1681685098
transform 1 0 128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_77
timestamp 1681685098
transform 1 0 136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_79
timestamp 1681685098
transform 1 0 144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_81
timestamp 1681685098
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_90
timestamp 1681685098
transform 1 0 160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_91
timestamp 1681685098
transform 1 0 168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_92
timestamp 1681685098
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use OR2X1  OR2X1_7
timestamp 1681685098
transform 1 0 184 0 -1 1770
box -8 -3 40 105
use XNOR2X1  XNOR2X1_6
timestamp 1681685098
transform -1 0 272 0 -1 1770
box -8 -3 64 105
use NAND3X1  NAND3X1_1
timestamp 1681685098
transform 1 0 272 0 -1 1770
box -8 -3 40 105
use FILL  FILL_93
timestamp 1681685098
transform 1 0 304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_94
timestamp 1681685098
transform 1 0 312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_96
timestamp 1681685098
transform 1 0 320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_98
timestamp 1681685098
transform 1 0 328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_103
timestamp 1681685098
transform 1 0 336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_104
timestamp 1681685098
transform 1 0 344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_105
timestamp 1681685098
transform 1 0 352 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_8
timestamp 1681685098
transform 1 0 360 0 -1 1770
box -8 -3 34 105
use FILL  FILL_106
timestamp 1681685098
transform 1 0 392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_107
timestamp 1681685098
transform 1 0 400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_108
timestamp 1681685098
transform 1 0 408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_109
timestamp 1681685098
transform 1 0 416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_110
timestamp 1681685098
transform 1 0 424 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1681685098
transform -1 0 464 0 -1 1770
box -8 -3 34 105
use INVX2  INVX2_9
timestamp 1681685098
transform -1 0 480 0 -1 1770
box -9 -3 26 105
use FILL  FILL_111
timestamp 1681685098
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_112
timestamp 1681685098
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_113
timestamp 1681685098
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_114
timestamp 1681685098
transform 1 0 504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_115
timestamp 1681685098
transform 1 0 512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_116
timestamp 1681685098
transform 1 0 520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_117
timestamp 1681685098
transform 1 0 528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_118
timestamp 1681685098
transform 1 0 536 0 -1 1770
box -8 -3 16 105
use OR2X1  OR2X1_9
timestamp 1681685098
transform 1 0 544 0 -1 1770
box -8 -3 40 105
use FILL  FILL_119
timestamp 1681685098
transform 1 0 576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_120
timestamp 1681685098
transform 1 0 584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_121
timestamp 1681685098
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_123
timestamp 1681685098
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_125
timestamp 1681685098
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_130
timestamp 1681685098
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1681685098
transform -1 0 656 0 -1 1770
box -8 -3 40 105
use INVX2  INVX2_11
timestamp 1681685098
transform -1 0 672 0 -1 1770
box -9 -3 26 105
use FILL  FILL_131
timestamp 1681685098
transform 1 0 672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_132
timestamp 1681685098
transform 1 0 680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_134
timestamp 1681685098
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_136
timestamp 1681685098
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use OR2X1  OR2X1_10
timestamp 1681685098
transform 1 0 704 0 -1 1770
box -8 -3 40 105
use XNOR2X1  XNOR2X1_8
timestamp 1681685098
transform 1 0 736 0 -1 1770
box -8 -3 64 105
use OAI21X1  OAI21X1_10
timestamp 1681685098
transform -1 0 824 0 -1 1770
box -8 -3 34 105
use FILL  FILL_149
timestamp 1681685098
transform 1 0 824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_154
timestamp 1681685098
transform 1 0 832 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_12
timestamp 1681685098
transform -1 0 856 0 -1 1770
box -9 -3 26 105
use FILL  FILL_155
timestamp 1681685098
transform 1 0 856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_157
timestamp 1681685098
transform 1 0 864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_162
timestamp 1681685098
transform 1 0 872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_163
timestamp 1681685098
transform 1 0 880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_164
timestamp 1681685098
transform 1 0 888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_165
timestamp 1681685098
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1681685098
transform 1 0 904 0 -1 1770
box -8 -3 32 105
use FILL  FILL_166
timestamp 1681685098
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_167
timestamp 1681685098
transform 1 0 936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_168
timestamp 1681685098
transform 1 0 944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_169
timestamp 1681685098
transform 1 0 952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_170
timestamp 1681685098
transform 1 0 960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_172
timestamp 1681685098
transform 1 0 968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_173
timestamp 1681685098
transform 1 0 976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_174
timestamp 1681685098
transform 1 0 984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_175
timestamp 1681685098
transform 1 0 992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_176
timestamp 1681685098
transform 1 0 1000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_177
timestamp 1681685098
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_12
timestamp 1681685098
transform -1 0 1048 0 -1 1770
box -8 -3 34 105
use INVX2  INVX2_13
timestamp 1681685098
transform 1 0 1048 0 -1 1770
box -9 -3 26 105
use FILL  FILL_178
timestamp 1681685098
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_179
timestamp 1681685098
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_180
timestamp 1681685098
transform 1 0 1080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_181
timestamp 1681685098
transform 1 0 1088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_182
timestamp 1681685098
transform 1 0 1096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_184
timestamp 1681685098
transform 1 0 1104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_186
timestamp 1681685098
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_192
timestamp 1681685098
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_2
timestamp 1681685098
transform -1 0 1152 0 -1 1770
box -8 -3 32 105
use FILL  FILL_193
timestamp 1681685098
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_194
timestamp 1681685098
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_195
timestamp 1681685098
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_196
timestamp 1681685098
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_198
timestamp 1681685098
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_3
timestamp 1681685098
transform 1 0 1192 0 -1 1770
box -8 -3 40 105
use FILL  FILL_202
timestamp 1681685098
transform 1 0 1224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_203
timestamp 1681685098
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_204
timestamp 1681685098
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_205
timestamp 1681685098
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_206
timestamp 1681685098
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_207
timestamp 1681685098
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_208
timestamp 1681685098
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_209
timestamp 1681685098
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_13
timestamp 1681685098
transform 1 0 1288 0 -1 1770
box -8 -3 34 105
use FILL  FILL_210
timestamp 1681685098
transform 1 0 1320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_211
timestamp 1681685098
transform 1 0 1328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_212
timestamp 1681685098
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_213
timestamp 1681685098
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_214
timestamp 1681685098
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_216
timestamp 1681685098
transform 1 0 1360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_218
timestamp 1681685098
transform 1 0 1368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_220
timestamp 1681685098
transform 1 0 1376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_252
timestamp 1681685098
transform 1 0 1384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_253
timestamp 1681685098
transform 1 0 1392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_254
timestamp 1681685098
transform 1 0 1400 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1681685098
transform 1 0 1408 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1681685098
transform 1 0 1504 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_16
timestamp 1681685098
transform -1 0 1616 0 -1 1770
box -9 -3 26 105
use XNOR2X1  XNOR2X1_9
timestamp 1681685098
transform 1 0 1616 0 -1 1770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_10
timestamp 1681685098
transform 1 0 1672 0 -1 1770
box -8 -3 64 105
use FILL  FILL_255
timestamp 1681685098
transform 1 0 1728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_256
timestamp 1681685098
transform 1 0 1736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_257
timestamp 1681685098
transform 1 0 1744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_258
timestamp 1681685098
transform 1 0 1752 0 -1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_6
timestamp 1681685098
transform 1 0 1760 0 -1 1770
box -8 -3 32 105
use FILL  FILL_260
timestamp 1681685098
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_262
timestamp 1681685098
transform 1 0 1792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_264
timestamp 1681685098
transform 1 0 1800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_266
timestamp 1681685098
transform 1 0 1808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_268
timestamp 1681685098
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_270
timestamp 1681685098
transform 1 0 1824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_272
timestamp 1681685098
transform 1 0 1832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_274
timestamp 1681685098
transform 1 0 1840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_275
timestamp 1681685098
transform 1 0 1848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_276
timestamp 1681685098
transform 1 0 1856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_277
timestamp 1681685098
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_15
timestamp 1681685098
transform -1 0 1904 0 -1 1770
box -8 -3 34 105
use FILL  FILL_278
timestamp 1681685098
transform 1 0 1904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_279
timestamp 1681685098
transform 1 0 1912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_280
timestamp 1681685098
transform 1 0 1920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_281
timestamp 1681685098
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_282
timestamp 1681685098
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_286
timestamp 1681685098
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1681685098
transform -1 0 1976 0 -1 1770
box -8 -3 32 105
use XNOR2X1  XNOR2X1_12
timestamp 1681685098
transform -1 0 2032 0 -1 1770
box -8 -3 64 105
use OR2X1  OR2X1_14
timestamp 1681685098
transform 1 0 2032 0 -1 1770
box -8 -3 40 105
use FILL  FILL_287
timestamp 1681685098
transform 1 0 2064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_289
timestamp 1681685098
transform 1 0 2072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_291
timestamp 1681685098
transform 1 0 2080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_293
timestamp 1681685098
transform 1 0 2088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_295
timestamp 1681685098
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_297
timestamp 1681685098
transform 1 0 2104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_299
timestamp 1681685098
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_301
timestamp 1681685098
transform 1 0 2120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_303
timestamp 1681685098
transform 1 0 2128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_305
timestamp 1681685098
transform 1 0 2136 0 -1 1770
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_7
timestamp 1681685098
transform 1 0 2194 0 1 1670
box -10 -3 10 3
use M2_M1  M2_M1_273
timestamp 1681685098
transform 1 0 132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1681685098
transform 1 0 132 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_187
timestamp 1681685098
transform 1 0 148 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_260
timestamp 1681685098
transform 1 0 148 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1681685098
transform 1 0 148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1681685098
transform 1 0 156 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_188
timestamp 1681685098
transform 1 0 212 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_261
timestamp 1681685098
transform 1 0 212 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_189
timestamp 1681685098
transform 1 0 244 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1681685098
transform 1 0 236 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1681685098
transform 1 0 268 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_275
timestamp 1681685098
transform 1 0 220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1681685098
transform 1 0 236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1681685098
transform 1 0 268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1681685098
transform 1 0 204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1681685098
transform 1 0 228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1681685098
transform 1 0 316 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_190
timestamp 1681685098
transform 1 0 332 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_262
timestamp 1681685098
transform 1 0 332 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1681685098
transform 1 0 380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1681685098
transform 1 0 372 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1681685098
transform 1 0 428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1681685098
transform 1 0 476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1681685098
transform 1 0 484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1681685098
transform 1 0 396 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1681685098
transform 1 0 484 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_191
timestamp 1681685098
transform 1 0 500 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_263
timestamp 1681685098
transform 1 0 500 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1681685098
transform 1 0 508 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_192
timestamp 1681685098
transform 1 0 540 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1681685098
transform 1 0 540 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_282
timestamp 1681685098
transform 1 0 564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1681685098
transform 1 0 580 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_216
timestamp 1681685098
transform 1 0 588 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1681685098
transform 1 0 620 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1681685098
transform 1 0 628 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_264
timestamp 1681685098
transform 1 0 628 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_194
timestamp 1681685098
transform 1 0 652 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_265
timestamp 1681685098
transform 1 0 660 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1681685098
transform 1 0 644 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1681685098
transform 1 0 652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1681685098
transform 1 0 628 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_217
timestamp 1681685098
transform 1 0 644 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1681685098
transform 1 0 660 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_316
timestamp 1681685098
transform 1 0 652 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_218
timestamp 1681685098
transform 1 0 652 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_266
timestamp 1681685098
transform 1 0 684 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1681685098
transform 1 0 708 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_219
timestamp 1681685098
transform 1 0 700 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1681685098
transform 1 0 836 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1681685098
transform 1 0 756 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1681685098
transform 1 0 860 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_285
timestamp 1681685098
transform 1 0 804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1681685098
transform 1 0 852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1681685098
transform 1 0 860 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1681685098
transform 1 0 756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1681685098
transform 1 0 772 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1681685098
transform 1 0 908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1681685098
transform 1 0 876 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1681685098
transform 1 0 892 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_220
timestamp 1681685098
transform 1 0 804 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1681685098
transform 1 0 820 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1681685098
transform 1 0 852 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1681685098
transform 1 0 892 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1681685098
transform 1 0 924 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1681685098
transform 1 0 948 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_322
timestamp 1681685098
transform 1 0 948 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1681685098
transform 1 0 964 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1681685098
transform 1 0 956 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1681685098
transform 1 0 996 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1681685098
transform 1 0 1020 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1681685098
transform 1 0 1052 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_289
timestamp 1681685098
transform 1 0 1004 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_195
timestamp 1681685098
transform 1 0 1028 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_323
timestamp 1681685098
transform 1 0 1020 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_237
timestamp 1681685098
transform 1 0 1044 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1681685098
transform 1 0 1076 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_324
timestamp 1681685098
transform 1 0 1076 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_203
timestamp 1681685098
transform 1 0 1228 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_290
timestamp 1681685098
transform 1 0 1188 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1681685098
transform 1 0 1220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1681685098
transform 1 0 1228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1681685098
transform 1 0 1140 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_196
timestamp 1681685098
transform 1 0 1292 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1681685098
transform 1 0 1284 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1681685098
transform 1 0 1252 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1681685098
transform 1 0 1268 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_293
timestamp 1681685098
transform 1 0 1284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1681685098
transform 1 0 1252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1681685098
transform 1 0 1260 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_224
timestamp 1681685098
transform 1 0 1252 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_328
timestamp 1681685098
transform 1 0 1316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1681685098
transform 1 0 1324 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_225
timestamp 1681685098
transform 1 0 1316 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1681685098
transform 1 0 1380 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_294
timestamp 1681685098
transform 1 0 1388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1681685098
transform 1 0 1380 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_183
timestamp 1681685098
transform 1 0 1412 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_268
timestamp 1681685098
transform 1 0 1404 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1681685098
transform 1 0 1412 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_212
timestamp 1681685098
transform 1 0 1420 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_270
timestamp 1681685098
transform 1 0 1492 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1681685098
transform 1 0 1468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1681685098
transform 1 0 1476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1681685098
transform 1 0 1460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1681685098
transform 1 0 1468 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_197
timestamp 1681685098
transform 1 0 1596 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1681685098
transform 1 0 1508 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_297
timestamp 1681685098
transform 1 0 1540 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_214
timestamp 1681685098
transform 1 0 1556 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_298
timestamp 1681685098
transform 1 0 1588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1681685098
transform 1 0 1596 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1681685098
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1681685098
transform 1 0 1492 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1681685098
transform 1 0 1508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1681685098
transform 1 0 1596 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_226
timestamp 1681685098
transform 1 0 1476 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1681685098
transform 1 0 1540 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1681685098
transform 1 0 1532 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1681685098
transform 1 0 1596 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1681685098
transform 1 0 1620 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_336
timestamp 1681685098
transform 1 0 1620 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_184
timestamp 1681685098
transform 1 0 1636 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_271
timestamp 1681685098
transform 1 0 1636 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1681685098
transform 1 0 1652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1681685098
transform 1 0 1716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1681685098
transform 1 0 1740 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_185
timestamp 1681685098
transform 1 0 1780 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_272
timestamp 1681685098
transform 1 0 1772 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1681685098
transform 1 0 1772 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_228
timestamp 1681685098
transform 1 0 1772 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1681685098
transform 1 0 1804 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_301
timestamp 1681685098
transform 1 0 1852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1681685098
transform 1 0 1900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1681685098
transform 1 0 1908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1681685098
transform 1 0 1820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1681685098
transform 1 0 1908 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_229
timestamp 1681685098
transform 1 0 1820 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1681685098
transform 1 0 1844 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1681685098
transform 1 0 1932 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_304
timestamp 1681685098
transform 1 0 2020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1681685098
transform 1 0 1980 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_232
timestamp 1681685098
transform 1 0 1980 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_346
timestamp 1681685098
transform 1 0 2084 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1681685098
transform 1 0 2124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1681685098
transform 1 0 2108 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_233
timestamp 1681685098
transform 1 0 2108 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1681685098
transform 1 0 2140 0 1 1595
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_8
timestamp 1681685098
transform 1 0 48 0 1 1570
box -10 -3 10 3
use FILL  FILL_306
timestamp 1681685098
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_307
timestamp 1681685098
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_308
timestamp 1681685098
transform 1 0 88 0 1 1570
box -8 -3 16 105
use FILL  FILL_309
timestamp 1681685098
transform 1 0 96 0 1 1570
box -8 -3 16 105
use FILL  FILL_310
timestamp 1681685098
transform 1 0 104 0 1 1570
box -8 -3 16 105
use FILL  FILL_311
timestamp 1681685098
transform 1 0 112 0 1 1570
box -8 -3 16 105
use FILL  FILL_312
timestamp 1681685098
transform 1 0 120 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_9
timestamp 1681685098
transform 1 0 128 0 1 1570
box -8 -3 32 105
use XNOR2X1  XNOR2X1_13
timestamp 1681685098
transform -1 0 208 0 1 1570
box -8 -3 64 105
use NAND2X1  NAND2X1_10
timestamp 1681685098
transform -1 0 232 0 1 1570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1681685098
transform -1 0 328 0 1 1570
box -8 -3 104 105
use FILL  FILL_313
timestamp 1681685098
transform 1 0 328 0 1 1570
box -8 -3 16 105
use FILL  FILL_327
timestamp 1681685098
transform 1 0 336 0 1 1570
box -8 -3 16 105
use FILL  FILL_329
timestamp 1681685098
transform 1 0 344 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_11
timestamp 1681685098
transform -1 0 376 0 1 1570
box -8 -3 32 105
use FILL  FILL_330
timestamp 1681685098
transform 1 0 376 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_240
timestamp 1681685098
transform 1 0 444 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1681685098
transform 1 0 476 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_15
timestamp 1681685098
transform 1 0 384 0 1 1570
box -8 -3 104 105
use M3_M2  M3_M2_242
timestamp 1681685098
transform 1 0 500 0 1 1575
box -3 -3 3 3
use NAND2X1  NAND2X1_12
timestamp 1681685098
transform 1 0 480 0 1 1570
box -8 -3 32 105
use FILL  FILL_331
timestamp 1681685098
transform 1 0 504 0 1 1570
box -8 -3 16 105
use FILL  FILL_338
timestamp 1681685098
transform 1 0 512 0 1 1570
box -8 -3 16 105
use FILL  FILL_340
timestamp 1681685098
transform 1 0 520 0 1 1570
box -8 -3 16 105
use FILL  FILL_341
timestamp 1681685098
transform 1 0 528 0 1 1570
box -8 -3 16 105
use FILL  FILL_342
timestamp 1681685098
transform 1 0 536 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_5
timestamp 1681685098
transform 1 0 544 0 1 1570
box -8 -3 32 105
use FILL  FILL_343
timestamp 1681685098
transform 1 0 568 0 1 1570
box -8 -3 16 105
use FILL  FILL_347
timestamp 1681685098
transform 1 0 576 0 1 1570
box -8 -3 16 105
use FILL  FILL_349
timestamp 1681685098
transform 1 0 584 0 1 1570
box -8 -3 16 105
use FILL  FILL_351
timestamp 1681685098
transform 1 0 592 0 1 1570
box -8 -3 16 105
use FILL  FILL_352
timestamp 1681685098
transform 1 0 600 0 1 1570
box -8 -3 16 105
use FILL  FILL_353
timestamp 1681685098
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_354
timestamp 1681685098
transform 1 0 616 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_17
timestamp 1681685098
transform -1 0 656 0 1 1570
box -8 -3 34 105
use FILL  FILL_355
timestamp 1681685098
transform 1 0 656 0 1 1570
box -8 -3 16 105
use FILL  FILL_356
timestamp 1681685098
transform 1 0 664 0 1 1570
box -8 -3 16 105
use FILL  FILL_357
timestamp 1681685098
transform 1 0 672 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_13
timestamp 1681685098
transform -1 0 704 0 1 1570
box -8 -3 32 105
use XNOR2X1  XNOR2X1_15
timestamp 1681685098
transform -1 0 760 0 1 1570
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1681685098
transform 1 0 760 0 1 1570
box -8 -3 104 105
use OR2X1  OR2X1_19
timestamp 1681685098
transform -1 0 888 0 1 1570
box -8 -3 40 105
use XNOR2X1  XNOR2X1_16
timestamp 1681685098
transform -1 0 944 0 1 1570
box -8 -3 64 105
use FILL  FILL_358
timestamp 1681685098
transform 1 0 944 0 1 1570
box -8 -3 16 105
use FILL  FILL_359
timestamp 1681685098
transform 1 0 952 0 1 1570
box -8 -3 16 105
use FILL  FILL_384
timestamp 1681685098
transform 1 0 960 0 1 1570
box -8 -3 16 105
use FILL  FILL_385
timestamp 1681685098
transform 1 0 968 0 1 1570
box -8 -3 16 105
use FILL  FILL_386
timestamp 1681685098
transform 1 0 976 0 1 1570
box -8 -3 16 105
use FILL  FILL_387
timestamp 1681685098
transform 1 0 984 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_14
timestamp 1681685098
transform -1 0 1016 0 1 1570
box -8 -3 32 105
use XNOR2X1  XNOR2X1_17
timestamp 1681685098
transform -1 0 1072 0 1 1570
box -8 -3 64 105
use FILL  FILL_388
timestamp 1681685098
transform 1 0 1072 0 1 1570
box -8 -3 16 105
use FILL  FILL_389
timestamp 1681685098
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_390
timestamp 1681685098
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use FILL  FILL_392
timestamp 1681685098
transform 1 0 1096 0 1 1570
box -8 -3 16 105
use FILL  FILL_394
timestamp 1681685098
transform 1 0 1104 0 1 1570
box -8 -3 16 105
use FILL  FILL_396
timestamp 1681685098
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_398
timestamp 1681685098
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_243
timestamp 1681685098
transform 1 0 1220 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_19
timestamp 1681685098
transform 1 0 1128 0 1 1570
box -8 -3 104 105
use FILL  FILL_400
timestamp 1681685098
transform 1 0 1224 0 1 1570
box -8 -3 16 105
use OR2X1  OR2X1_20
timestamp 1681685098
transform -1 0 1264 0 1 1570
box -8 -3 40 105
use M3_M2  M3_M2_244
timestamp 1681685098
transform 1 0 1324 0 1 1575
box -3 -3 3 3
use XNOR2X1  XNOR2X1_18
timestamp 1681685098
transform -1 0 1320 0 1 1570
box -8 -3 64 105
use INVX2  INVX2_18
timestamp 1681685098
transform 1 0 1320 0 1 1570
box -9 -3 26 105
use FILL  FILL_401
timestamp 1681685098
transform 1 0 1336 0 1 1570
box -8 -3 16 105
use FILL  FILL_402
timestamp 1681685098
transform 1 0 1344 0 1 1570
box -8 -3 16 105
use FILL  FILL_403
timestamp 1681685098
transform 1 0 1352 0 1 1570
box -8 -3 16 105
use FILL  FILL_420
timestamp 1681685098
transform 1 0 1360 0 1 1570
box -8 -3 16 105
use FILL  FILL_422
timestamp 1681685098
transform 1 0 1368 0 1 1570
box -8 -3 16 105
use FILL  FILL_424
timestamp 1681685098
transform 1 0 1376 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_15
timestamp 1681685098
transform 1 0 1384 0 1 1570
box -8 -3 32 105
use FILL  FILL_426
timestamp 1681685098
transform 1 0 1408 0 1 1570
box -8 -3 16 105
use FILL  FILL_429
timestamp 1681685098
transform 1 0 1416 0 1 1570
box -8 -3 16 105
use FILL  FILL_431
timestamp 1681685098
transform 1 0 1424 0 1 1570
box -8 -3 16 105
use FILL  FILL_433
timestamp 1681685098
transform 1 0 1432 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_16
timestamp 1681685098
transform -1 0 1464 0 1 1570
box -8 -3 32 105
use OAI21X1  OAI21X1_21
timestamp 1681685098
transform 1 0 1464 0 1 1570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1681685098
transform 1 0 1496 0 1 1570
box -8 -3 104 105
use OAI21X1  OAI21X1_22
timestamp 1681685098
transform 1 0 1592 0 1 1570
box -8 -3 34 105
use FILL  FILL_434
timestamp 1681685098
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_17
timestamp 1681685098
transform -1 0 1656 0 1 1570
box -8 -3 32 105
use FILL  FILL_435
timestamp 1681685098
transform 1 0 1656 0 1 1570
box -8 -3 16 105
use FILL  FILL_436
timestamp 1681685098
transform 1 0 1664 0 1 1570
box -8 -3 16 105
use FILL  FILL_437
timestamp 1681685098
transform 1 0 1672 0 1 1570
box -8 -3 16 105
use FILL  FILL_438
timestamp 1681685098
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use FILL  FILL_439
timestamp 1681685098
transform 1 0 1688 0 1 1570
box -8 -3 16 105
use FILL  FILL_440
timestamp 1681685098
transform 1 0 1696 0 1 1570
box -8 -3 16 105
use FILL  FILL_441
timestamp 1681685098
transform 1 0 1704 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_21
timestamp 1681685098
transform 1 0 1712 0 1 1570
box -9 -3 26 105
use FILL  FILL_442
timestamp 1681685098
transform 1 0 1728 0 1 1570
box -8 -3 16 105
use FILL  FILL_443
timestamp 1681685098
transform 1 0 1736 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_23
timestamp 1681685098
transform 1 0 1744 0 1 1570
box -8 -3 34 105
use FILL  FILL_444
timestamp 1681685098
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use FILL  FILL_445
timestamp 1681685098
transform 1 0 1784 0 1 1570
box -8 -3 16 105
use FILL  FILL_446
timestamp 1681685098
transform 1 0 1792 0 1 1570
box -8 -3 16 105
use FILL  FILL_447
timestamp 1681685098
transform 1 0 1800 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1681685098
transform 1 0 1808 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_22
timestamp 1681685098
transform 1 0 1904 0 1 1570
box -9 -3 26 105
use FILL  FILL_448
timestamp 1681685098
transform 1 0 1920 0 1 1570
box -8 -3 16 105
use FILL  FILL_449
timestamp 1681685098
transform 1 0 1928 0 1 1570
box -8 -3 16 105
use FILL  FILL_480
timestamp 1681685098
transform 1 0 1936 0 1 1570
box -8 -3 16 105
use FILL  FILL_482
timestamp 1681685098
transform 1 0 1944 0 1 1570
box -8 -3 16 105
use FILL  FILL_484
timestamp 1681685098
transform 1 0 1952 0 1 1570
box -8 -3 16 105
use FILL  FILL_485
timestamp 1681685098
transform 1 0 1960 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1681685098
transform 1 0 1968 0 1 1570
box -8 -3 104 105
use FILL  FILL_486
timestamp 1681685098
transform 1 0 2064 0 1 1570
box -8 -3 16 105
use FILL  FILL_489
timestamp 1681685098
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_490
timestamp 1681685098
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_491
timestamp 1681685098
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use OR2X1  OR2X1_22
timestamp 1681685098
transform 1 0 2096 0 1 1570
box -8 -3 40 105
use FILL  FILL_492
timestamp 1681685098
transform 1 0 2128 0 1 1570
box -8 -3 16 105
use FILL  FILL_493
timestamp 1681685098
transform 1 0 2136 0 1 1570
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_9
timestamp 1681685098
transform 1 0 2170 0 1 1570
box -10 -3 10 3
use M3_M2  M3_M2_250
timestamp 1681685098
transform 1 0 84 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_347
timestamp 1681685098
transform 1 0 172 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1681685098
transform 1 0 84 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1681685098
transform 1 0 180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1681685098
transform 1 0 116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1681685098
transform 1 0 164 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_283
timestamp 1681685098
transform 1 0 180 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_421
timestamp 1681685098
transform 1 0 220 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_284
timestamp 1681685098
transform 1 0 220 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_388
timestamp 1681685098
transform 1 0 252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1681685098
transform 1 0 260 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1681685098
transform 1 0 284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1681685098
transform 1 0 284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1681685098
transform 1 0 348 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_285
timestamp 1681685098
transform 1 0 348 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_348
timestamp 1681685098
transform 1 0 380 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_251
timestamp 1681685098
transform 1 0 396 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_391
timestamp 1681685098
transform 1 0 404 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_245
timestamp 1681685098
transform 1 0 484 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1681685098
transform 1 0 436 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_349
timestamp 1681685098
transform 1 0 444 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_253
timestamp 1681685098
transform 1 0 452 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_358
timestamp 1681685098
transform 1 0 452 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_286
timestamp 1681685098
transform 1 0 444 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1681685098
transform 1 0 508 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_359
timestamp 1681685098
transform 1 0 500 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1681685098
transform 1 0 500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1681685098
transform 1 0 508 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_275
timestamp 1681685098
transform 1 0 500 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1681685098
transform 1 0 524 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_360
timestamp 1681685098
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_266
timestamp 1681685098
transform 1 0 532 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1681685098
transform 1 0 524 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_350
timestamp 1681685098
transform 1 0 564 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_267
timestamp 1681685098
transform 1 0 564 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_361
timestamp 1681685098
transform 1 0 604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1681685098
transform 1 0 628 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_287
timestamp 1681685098
transform 1 0 604 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_362
timestamp 1681685098
transform 1 0 700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1681685098
transform 1 0 692 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1681685098
transform 1 0 700 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_288
timestamp 1681685098
transform 1 0 732 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_363
timestamp 1681685098
transform 1 0 756 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_289
timestamp 1681685098
transform 1 0 772 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1681685098
transform 1 0 844 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_422
timestamp 1681685098
transform 1 0 828 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1681685098
transform 1 0 836 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1681685098
transform 1 0 892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1681685098
transform 1 0 900 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_294
timestamp 1681685098
transform 1 0 900 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_398
timestamp 1681685098
transform 1 0 916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1681685098
transform 1 0 940 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1681685098
transform 1 0 932 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1681685098
transform 1 0 948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1681685098
transform 1 0 964 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_255
timestamp 1681685098
transform 1 0 988 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1681685098
transform 1 0 1028 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1681685098
transform 1 0 1076 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_366
timestamp 1681685098
transform 1 0 988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1681685098
transform 1 0 1076 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1681685098
transform 1 0 996 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1681685098
transform 1 0 1028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1681685098
transform 1 0 988 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_258
timestamp 1681685098
transform 1 0 1140 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_368
timestamp 1681685098
transform 1 0 1132 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_290
timestamp 1681685098
transform 1 0 1132 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_402
timestamp 1681685098
transform 1 0 1156 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1681685098
transform 1 0 1188 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1681685098
transform 1 0 1220 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1681685098
transform 1 0 1244 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_277
timestamp 1681685098
transform 1 0 1244 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1681685098
transform 1 0 1268 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1681685098
transform 1 0 1276 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_404
timestamp 1681685098
transform 1 0 1308 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_269
timestamp 1681685098
transform 1 0 1316 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_405
timestamp 1681685098
transform 1 0 1324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1681685098
transform 1 0 1316 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1681685098
transform 1 0 1300 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_295
timestamp 1681685098
transform 1 0 1300 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1681685098
transform 1 0 1324 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_351
timestamp 1681685098
transform 1 0 1348 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1681685098
transform 1 0 1372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1681685098
transform 1 0 1380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1681685098
transform 1 0 1364 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_296
timestamp 1681685098
transform 1 0 1364 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_372
timestamp 1681685098
transform 1 0 1396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1681685098
transform 1 0 1452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1681685098
transform 1 0 1468 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_270
timestamp 1681685098
transform 1 0 1460 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_407
timestamp 1681685098
transform 1 0 1468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1681685098
transform 1 0 1484 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_279
timestamp 1681685098
transform 1 0 1484 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_375
timestamp 1681685098
transform 1 0 1508 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_271
timestamp 1681685098
transform 1 0 1500 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_409
timestamp 1681685098
transform 1 0 1508 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_280
timestamp 1681685098
transform 1 0 1508 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1681685098
transform 1 0 1596 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_376
timestamp 1681685098
transform 1 0 1596 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_247
timestamp 1681685098
transform 1 0 1692 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1681685098
transform 1 0 1740 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1681685098
transform 1 0 1732 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_377
timestamp 1681685098
transform 1 0 1732 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1681685098
transform 1 0 1652 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1681685098
transform 1 0 1700 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_272
timestamp 1681685098
transform 1 0 1732 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_352
timestamp 1681685098
transform 1 0 1748 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_263
timestamp 1681685098
transform 1 0 1748 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1681685098
transform 1 0 1820 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_378
timestamp 1681685098
transform 1 0 1804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1681685098
transform 1 0 1788 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1681685098
transform 1 0 1812 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1681685098
transform 1 0 1820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1681685098
transform 1 0 1852 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_281
timestamp 1681685098
transform 1 0 1812 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1681685098
transform 1 0 1852 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1681685098
transform 1 0 1804 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1681685098
transform 1 0 1820 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_379
timestamp 1681685098
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1681685098
transform 1 0 1900 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1681685098
transform 1 0 1900 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_298
timestamp 1681685098
transform 1 0 1900 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_428
timestamp 1681685098
transform 1 0 1940 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1681685098
transform 1 0 1956 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_249
timestamp 1681685098
transform 1 0 1996 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1681685098
transform 1 0 1988 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_381
timestamp 1681685098
transform 1 0 1996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1681685098
transform 1 0 2020 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1681685098
transform 1 0 1980 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1681685098
transform 1 0 1996 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_273
timestamp 1681685098
transform 1 0 2004 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_429
timestamp 1681685098
transform 1 0 1988 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1681685098
transform 1 0 1972 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1681685098
transform 1 0 2044 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_265
timestamp 1681685098
transform 1 0 2052 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1681685098
transform 1 0 2036 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_419
timestamp 1681685098
transform 1 0 2052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1681685098
transform 1 0 2060 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1681685098
transform 1 0 2028 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_293
timestamp 1681685098
transform 1 0 2028 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_384
timestamp 1681685098
transform 1 0 2084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1681685098
transform 1 0 2140 0 1 1535
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_10
timestamp 1681685098
transform 1 0 24 0 1 1470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_14
timestamp 1681685098
transform 1 0 72 0 -1 1570
box -8 -3 104 105
use OR2X1  OR2X1_15
timestamp 1681685098
transform 1 0 168 0 -1 1570
box -8 -3 40 105
use FILL  FILL_314
timestamp 1681685098
transform 1 0 200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_315
timestamp 1681685098
transform 1 0 208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_316
timestamp 1681685098
transform 1 0 216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_317
timestamp 1681685098
transform 1 0 224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_318
timestamp 1681685098
transform 1 0 232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_319
timestamp 1681685098
transform 1 0 240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_320
timestamp 1681685098
transform 1 0 248 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_16
timestamp 1681685098
transform -1 0 288 0 -1 1570
box -8 -3 34 105
use FILL  FILL_321
timestamp 1681685098
transform 1 0 288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_322
timestamp 1681685098
transform 1 0 296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_323
timestamp 1681685098
transform 1 0 304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_324
timestamp 1681685098
transform 1 0 312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_325
timestamp 1681685098
transform 1 0 320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_326
timestamp 1681685098
transform 1 0 328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_328
timestamp 1681685098
transform 1 0 336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_332
timestamp 1681685098
transform 1 0 344 0 -1 1570
box -8 -3 16 105
use OR2X1  OR2X1_16
timestamp 1681685098
transform -1 0 384 0 -1 1570
box -8 -3 40 105
use FILL  FILL_333
timestamp 1681685098
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_334
timestamp 1681685098
transform 1 0 392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_335
timestamp 1681685098
transform 1 0 400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_336
timestamp 1681685098
transform 1 0 408 0 -1 1570
box -8 -3 16 105
use OR2X1  OR2X1_17
timestamp 1681685098
transform -1 0 448 0 -1 1570
box -8 -3 40 105
use XNOR2X1  XNOR2X1_14
timestamp 1681685098
transform 1 0 448 0 -1 1570
box -8 -3 64 105
use FILL  FILL_337
timestamp 1681685098
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_339
timestamp 1681685098
transform 1 0 512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_344
timestamp 1681685098
transform 1 0 520 0 -1 1570
box -8 -3 16 105
use OR2X1  OR2X1_18
timestamp 1681685098
transform -1 0 560 0 -1 1570
box -8 -3 40 105
use FILL  FILL_345
timestamp 1681685098
transform 1 0 560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_346
timestamp 1681685098
transform 1 0 568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_348
timestamp 1681685098
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_350
timestamp 1681685098
transform 1 0 584 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1681685098
transform 1 0 592 0 -1 1570
box -8 -3 104 105
use FILL  FILL_360
timestamp 1681685098
transform 1 0 688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_361
timestamp 1681685098
transform 1 0 696 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_18
timestamp 1681685098
transform 1 0 704 0 -1 1570
box -8 -3 34 105
use FILL  FILL_362
timestamp 1681685098
transform 1 0 736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_363
timestamp 1681685098
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_364
timestamp 1681685098
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_365
timestamp 1681685098
transform 1 0 760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_366
timestamp 1681685098
transform 1 0 768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_367
timestamp 1681685098
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_368
timestamp 1681685098
transform 1 0 784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_369
timestamp 1681685098
transform 1 0 792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_370
timestamp 1681685098
transform 1 0 800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_371
timestamp 1681685098
transform 1 0 808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_372
timestamp 1681685098
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_373
timestamp 1681685098
transform 1 0 824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_374
timestamp 1681685098
transform 1 0 832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_375
timestamp 1681685098
transform 1 0 840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_376
timestamp 1681685098
transform 1 0 848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_377
timestamp 1681685098
transform 1 0 856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_378
timestamp 1681685098
transform 1 0 864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_379
timestamp 1681685098
transform 1 0 872 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1681685098
transform 1 0 880 0 -1 1570
box -8 -3 40 105
use FILL  FILL_380
timestamp 1681685098
transform 1 0 912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_381
timestamp 1681685098
transform 1 0 920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_382
timestamp 1681685098
transform 1 0 928 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_17
timestamp 1681685098
transform 1 0 936 0 -1 1570
box -9 -3 26 105
use FILL  FILL_383
timestamp 1681685098
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_19
timestamp 1681685098
transform 1 0 960 0 -1 1570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1681685098
transform -1 0 1088 0 -1 1570
box -8 -3 104 105
use FILL  FILL_391
timestamp 1681685098
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_393
timestamp 1681685098
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_395
timestamp 1681685098
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_397
timestamp 1681685098
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_399
timestamp 1681685098
transform 1 0 1120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_404
timestamp 1681685098
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_19
timestamp 1681685098
transform 1 0 1136 0 -1 1570
box -9 -3 26 105
use FILL  FILL_405
timestamp 1681685098
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_406
timestamp 1681685098
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_407
timestamp 1681685098
transform 1 0 1168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_408
timestamp 1681685098
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_409
timestamp 1681685098
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_410
timestamp 1681685098
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_411
timestamp 1681685098
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_412
timestamp 1681685098
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_413
timestamp 1681685098
transform 1 0 1216 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_20
timestamp 1681685098
transform -1 0 1256 0 -1 1570
box -8 -3 34 105
use FILL  FILL_414
timestamp 1681685098
transform 1 0 1256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_415
timestamp 1681685098
transform 1 0 1264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_416
timestamp 1681685098
transform 1 0 1272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_417
timestamp 1681685098
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_5
timestamp 1681685098
transform -1 0 1320 0 -1 1570
box -8 -3 40 105
use FILL  FILL_418
timestamp 1681685098
transform 1 0 1320 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_6
timestamp 1681685098
transform -1 0 1352 0 -1 1570
box -8 -3 32 105
use FILL  FILL_419
timestamp 1681685098
transform 1 0 1352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_421
timestamp 1681685098
transform 1 0 1360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_423
timestamp 1681685098
transform 1 0 1368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_425
timestamp 1681685098
transform 1 0 1376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_427
timestamp 1681685098
transform 1 0 1384 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_20
timestamp 1681685098
transform 1 0 1392 0 -1 1570
box -9 -3 26 105
use FILL  FILL_428
timestamp 1681685098
transform 1 0 1408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_430
timestamp 1681685098
transform 1 0 1416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_432
timestamp 1681685098
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_450
timestamp 1681685098
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_451
timestamp 1681685098
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_452
timestamp 1681685098
transform 1 0 1448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_453
timestamp 1681685098
transform 1 0 1456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_454
timestamp 1681685098
transform 1 0 1464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_455
timestamp 1681685098
transform 1 0 1472 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_0
timestamp 1681685098
transform 1 0 1480 0 -1 1570
box -5 -3 28 105
use FILL  FILL_456
timestamp 1681685098
transform 1 0 1504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_457
timestamp 1681685098
transform 1 0 1512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_458
timestamp 1681685098
transform 1 0 1520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_459
timestamp 1681685098
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_460
timestamp 1681685098
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_461
timestamp 1681685098
transform 1 0 1544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_462
timestamp 1681685098
transform 1 0 1552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_463
timestamp 1681685098
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_464
timestamp 1681685098
transform 1 0 1568 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_1
timestamp 1681685098
transform 1 0 1576 0 -1 1570
box -5 -3 28 105
use FILL  FILL_465
timestamp 1681685098
transform 1 0 1600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_466
timestamp 1681685098
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_467
timestamp 1681685098
transform 1 0 1616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_468
timestamp 1681685098
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_469
timestamp 1681685098
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_470
timestamp 1681685098
transform 1 0 1640 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1681685098
transform -1 0 1744 0 -1 1570
box -8 -3 104 105
use FILL  FILL_471
timestamp 1681685098
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_472
timestamp 1681685098
transform 1 0 1752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_473
timestamp 1681685098
transform 1 0 1760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_474
timestamp 1681685098
transform 1 0 1768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_475
timestamp 1681685098
transform 1 0 1776 0 -1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_2
timestamp 1681685098
transform -1 0 1816 0 -1 1570
box -7 -3 39 105
use XNOR2X1  XNOR2X1_19
timestamp 1681685098
transform 1 0 1816 0 -1 1570
box -8 -3 64 105
use FILL  FILL_476
timestamp 1681685098
transform 1 0 1872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_477
timestamp 1681685098
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_478
timestamp 1681685098
transform 1 0 1888 0 -1 1570
box -8 -3 16 105
use OR2X1  OR2X1_21
timestamp 1681685098
transform 1 0 1896 0 -1 1570
box -8 -3 40 105
use FILL  FILL_479
timestamp 1681685098
transform 1 0 1928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_481
timestamp 1681685098
transform 1 0 1936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_483
timestamp 1681685098
transform 1 0 1944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_487
timestamp 1681685098
transform 1 0 1952 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_6
timestamp 1681685098
transform -1 0 1992 0 -1 1570
box -8 -3 40 105
use OAI21X1  OAI21X1_24
timestamp 1681685098
transform 1 0 1992 0 -1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_18
timestamp 1681685098
transform -1 0 2048 0 -1 1570
box -8 -3 32 105
use INVX2  INVX2_23
timestamp 1681685098
transform -1 0 2064 0 -1 1570
box -9 -3 26 105
use FILL  FILL_488
timestamp 1681685098
transform 1 0 2064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_494
timestamp 1681685098
transform 1 0 2072 0 -1 1570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_20
timestamp 1681685098
transform -1 0 2136 0 -1 1570
box -8 -3 64 105
use FILL  FILL_495
timestamp 1681685098
transform 1 0 2136 0 -1 1570
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_11
timestamp 1681685098
transform 1 0 2194 0 1 1470
box -10 -3 10 3
use M3_M2  M3_M2_306
timestamp 1681685098
transform 1 0 244 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1681685098
transform 1 0 236 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_436
timestamp 1681685098
transform 1 0 244 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1681685098
transform 1 0 132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1681685098
transform 1 0 172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1681685098
transform 1 0 188 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_324
timestamp 1681685098
transform 1 0 196 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1681685098
transform 1 0 228 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_456
timestamp 1681685098
transform 1 0 236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1681685098
transform 1 0 84 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1681685098
transform 1 0 172 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_340
timestamp 1681685098
transform 1 0 132 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_485
timestamp 1681685098
transform 1 0 220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1681685098
transform 1 0 228 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_341
timestamp 1681685098
transform 1 0 220 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1681685098
transform 1 0 260 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_487
timestamp 1681685098
transform 1 0 260 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1681685098
transform 1 0 284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1681685098
transform 1 0 340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1681685098
transform 1 0 372 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_326
timestamp 1681685098
transform 1 0 380 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_459
timestamp 1681685098
transform 1 0 404 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_327
timestamp 1681685098
transform 1 0 412 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1681685098
transform 1 0 428 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_437
timestamp 1681685098
transform 1 0 428 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1681685098
transform 1 0 420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1681685098
transform 1 0 356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1681685098
transform 1 0 412 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_350
timestamp 1681685098
transform 1 0 388 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1681685098
transform 1 0 420 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_438
timestamp 1681685098
transform 1 0 452 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_328
timestamp 1681685098
transform 1 0 452 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1681685098
transform 1 0 484 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_491
timestamp 1681685098
transform 1 0 484 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_309
timestamp 1681685098
transform 1 0 548 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_439
timestamp 1681685098
transform 1 0 556 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1681685098
transform 1 0 548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1681685098
transform 1 0 532 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_329
timestamp 1681685098
transform 1 0 556 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_493
timestamp 1681685098
transform 1 0 628 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_310
timestamp 1681685098
transform 1 0 660 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_462
timestamp 1681685098
transform 1 0 700 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1681685098
transform 1 0 708 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_352
timestamp 1681685098
transform 1 0 708 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_440
timestamp 1681685098
transform 1 0 836 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1681685098
transform 1 0 756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1681685098
transform 1 0 812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1681685098
transform 1 0 828 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1681685098
transform 1 0 732 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1681685098
transform 1 0 820 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_342
timestamp 1681685098
transform 1 0 732 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1681685098
transform 1 0 836 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1681685098
transform 1 0 812 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1681685098
transform 1 0 828 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1681685098
transform 1 0 940 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1681685098
transform 1 0 884 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_466
timestamp 1681685098
transform 1 0 908 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1681685098
transform 1 0 940 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1681685098
transform 1 0 956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1681685098
transform 1 0 860 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1681685098
transform 1 0 948 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_343
timestamp 1681685098
transform 1 0 860 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1681685098
transform 1 0 908 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_499
timestamp 1681685098
transform 1 0 972 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_345
timestamp 1681685098
transform 1 0 972 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_469
timestamp 1681685098
transform 1 0 988 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_355
timestamp 1681685098
transform 1 0 980 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_500
timestamp 1681685098
transform 1 0 996 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_304
timestamp 1681685098
transform 1 0 1036 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1681685098
transform 1 0 1028 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1681685098
transform 1 0 1052 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_441
timestamp 1681685098
transform 1 0 1012 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1681685098
transform 1 0 1028 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1681685098
transform 1 0 1036 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_332
timestamp 1681685098
transform 1 0 1012 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1681685098
transform 1 0 1028 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_470
timestamp 1681685098
transform 1 0 1052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1681685098
transform 1 0 1028 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_305
timestamp 1681685098
transform 1 0 1084 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1681685098
transform 1 0 1076 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_471
timestamp 1681685098
transform 1 0 1068 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1681685098
transform 1 0 1060 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1681685098
transform 1 0 1092 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_356
timestamp 1681685098
transform 1 0 1092 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_504
timestamp 1681685098
transform 1 0 1140 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1681685098
transform 1 0 1164 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1681685098
transform 1 0 1180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1681685098
transform 1 0 1212 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1681685098
transform 1 0 1220 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_314
timestamp 1681685098
transform 1 0 1252 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_472
timestamp 1681685098
transform 1 0 1252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1681685098
transform 1 0 1268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1681685098
transform 1 0 1284 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1681685098
transform 1 0 1348 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_315
timestamp 1681685098
transform 1 0 1380 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_447
timestamp 1681685098
transform 1 0 1396 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1681685098
transform 1 0 1412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1681685098
transform 1 0 1428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1681685098
transform 1 0 1412 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1681685098
transform 1 0 1468 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1681685098
transform 1 0 1476 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_334
timestamp 1681685098
transform 1 0 1476 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_510
timestamp 1681685098
transform 1 0 1468 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_320
timestamp 1681685098
transform 1 0 1492 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1681685098
transform 1 0 1532 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_475
timestamp 1681685098
transform 1 0 1500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1681685098
transform 1 0 1532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1681685098
transform 1 0 1580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1681685098
transform 1 0 1652 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_346
timestamp 1681685098
transform 1 0 1652 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_477
timestamp 1681685098
transform 1 0 1684 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_335
timestamp 1681685098
transform 1 0 1692 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_513
timestamp 1681685098
transform 1 0 1676 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1681685098
transform 1 0 1700 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_347
timestamp 1681685098
transform 1 0 1684 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_449
timestamp 1681685098
transform 1 0 1708 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1681685098
transform 1 0 1716 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_336
timestamp 1681685098
transform 1 0 1716 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_435
timestamp 1681685098
transform 1 0 1804 0 1 1435
box -2 -2 2 2
use M3_M2  M3_M2_316
timestamp 1681685098
transform 1 0 1812 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1681685098
transform 1 0 1836 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1681685098
transform 1 0 1804 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_451
timestamp 1681685098
transform 1 0 1812 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_337
timestamp 1681685098
transform 1 0 1812 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_478
timestamp 1681685098
transform 1 0 1820 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1681685098
transform 1 0 1796 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_323
timestamp 1681685098
transform 1 0 1844 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_516
timestamp 1681685098
transform 1 0 1836 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1681685098
transform 1 0 1844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1681685098
transform 1 0 1884 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_299
timestamp 1681685098
transform 1 0 1900 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_521
timestamp 1681685098
transform 1 0 1900 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_300
timestamp 1681685098
transform 1 0 1940 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1681685098
transform 1 0 1988 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1681685098
transform 1 0 2028 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_480
timestamp 1681685098
transform 1 0 1980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1681685098
transform 1 0 2012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1681685098
transform 1 0 2028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1681685098
transform 1 0 1932 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_338
timestamp 1681685098
transform 1 0 1980 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_522
timestamp 1681685098
transform 1 0 1916 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1681685098
transform 1 0 2036 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_339
timestamp 1681685098
transform 1 0 2052 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_520
timestamp 1681685098
transform 1 0 2060 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_348
timestamp 1681685098
transform 1 0 2028 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_452
timestamp 1681685098
transform 1 0 2068 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_349
timestamp 1681685098
transform 1 0 2068 0 1 1395
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_12
timestamp 1681685098
transform 1 0 48 0 1 1370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_24
timestamp 1681685098
transform 1 0 72 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_357
timestamp 1681685098
transform 1 0 196 0 1 1375
box -3 -3 3 3
use XNOR2X1  XNOR2X1_21
timestamp 1681685098
transform -1 0 224 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_358
timestamp 1681685098
transform 1 0 252 0 1 1375
box -3 -3 3 3
use NAND2X1  NAND2X1_19
timestamp 1681685098
transform 1 0 224 0 1 1370
box -8 -3 32 105
use FILL  FILL_496
timestamp 1681685098
transform 1 0 248 0 1 1370
box -8 -3 16 105
use FILL  FILL_498
timestamp 1681685098
transform 1 0 256 0 1 1370
box -8 -3 16 105
use FILL  FILL_500
timestamp 1681685098
transform 1 0 264 0 1 1370
box -8 -3 16 105
use FILL  FILL_502
timestamp 1681685098
transform 1 0 272 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_25
timestamp 1681685098
transform 1 0 280 0 1 1370
box -9 -3 26 105
use FILL  FILL_503
timestamp 1681685098
transform 1 0 296 0 1 1370
box -8 -3 16 105
use FILL  FILL_504
timestamp 1681685098
transform 1 0 304 0 1 1370
box -8 -3 16 105
use FILL  FILL_507
timestamp 1681685098
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_509
timestamp 1681685098
transform 1 0 320 0 1 1370
box -8 -3 16 105
use FILL  FILL_510
timestamp 1681685098
transform 1 0 328 0 1 1370
box -8 -3 16 105
use FILL  FILL_511
timestamp 1681685098
transform 1 0 336 0 1 1370
box -8 -3 16 105
use FILL  FILL_512
timestamp 1681685098
transform 1 0 344 0 1 1370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_22
timestamp 1681685098
transform -1 0 408 0 1 1370
box -8 -3 64 105
use NAND2X1  NAND2X1_20
timestamp 1681685098
transform 1 0 408 0 1 1370
box -8 -3 32 105
use FILL  FILL_513
timestamp 1681685098
transform 1 0 432 0 1 1370
box -8 -3 16 105
use FILL  FILL_514
timestamp 1681685098
transform 1 0 440 0 1 1370
box -8 -3 16 105
use FILL  FILL_515
timestamp 1681685098
transform 1 0 448 0 1 1370
box -8 -3 16 105
use FILL  FILL_516
timestamp 1681685098
transform 1 0 456 0 1 1370
box -8 -3 16 105
use FILL  FILL_517
timestamp 1681685098
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_518
timestamp 1681685098
transform 1 0 472 0 1 1370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_23
timestamp 1681685098
transform 1 0 480 0 1 1370
box -8 -3 64 105
use NAND2X1  NAND2X1_21
timestamp 1681685098
transform 1 0 536 0 1 1370
box -8 -3 32 105
use FILL  FILL_519
timestamp 1681685098
transform 1 0 560 0 1 1370
box -8 -3 16 105
use FILL  FILL_520
timestamp 1681685098
transform 1 0 568 0 1 1370
box -8 -3 16 105
use FILL  FILL_521
timestamp 1681685098
transform 1 0 576 0 1 1370
box -8 -3 16 105
use FILL  FILL_527
timestamp 1681685098
transform 1 0 584 0 1 1370
box -8 -3 16 105
use FILL  FILL_529
timestamp 1681685098
transform 1 0 592 0 1 1370
box -8 -3 16 105
use FILL  FILL_531
timestamp 1681685098
transform 1 0 600 0 1 1370
box -8 -3 16 105
use FILL  FILL_532
timestamp 1681685098
transform 1 0 608 0 1 1370
box -8 -3 16 105
use FILL  FILL_533
timestamp 1681685098
transform 1 0 616 0 1 1370
box -8 -3 16 105
use FILL  FILL_534
timestamp 1681685098
transform 1 0 624 0 1 1370
box -8 -3 16 105
use FILL  FILL_535
timestamp 1681685098
transform 1 0 632 0 1 1370
box -8 -3 16 105
use FILL  FILL_536
timestamp 1681685098
transform 1 0 640 0 1 1370
box -8 -3 16 105
use FILL  FILL_539
timestamp 1681685098
transform 1 0 648 0 1 1370
box -8 -3 16 105
use FILL  FILL_541
timestamp 1681685098
transform 1 0 656 0 1 1370
box -8 -3 16 105
use FILL  FILL_543
timestamp 1681685098
transform 1 0 664 0 1 1370
box -8 -3 16 105
use FILL  FILL_544
timestamp 1681685098
transform 1 0 672 0 1 1370
box -8 -3 16 105
use FILL  FILL_545
timestamp 1681685098
transform 1 0 680 0 1 1370
box -8 -3 16 105
use FILL  FILL_546
timestamp 1681685098
transform 1 0 688 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_28
timestamp 1681685098
transform -1 0 712 0 1 1370
box -9 -3 26 105
use FILL  FILL_547
timestamp 1681685098
transform 1 0 712 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1681685098
transform 1 0 720 0 1 1370
box -8 -3 104 105
use NAND2X1  NAND2X1_22
timestamp 1681685098
transform 1 0 816 0 1 1370
box -8 -3 32 105
use FILL  FILL_548
timestamp 1681685098
transform 1 0 840 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1681685098
transform 1 0 848 0 1 1370
box -8 -3 104 105
use OAI21X1  OAI21X1_28
timestamp 1681685098
transform 1 0 944 0 1 1370
box -8 -3 34 105
use FILL  FILL_555
timestamp 1681685098
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_566
timestamp 1681685098
transform 1 0 984 0 1 1370
box -8 -3 16 105
use FILL  FILL_568
timestamp 1681685098
transform 1 0 992 0 1 1370
box -8 -3 16 105
use FILL  FILL_570
timestamp 1681685098
transform 1 0 1000 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_24
timestamp 1681685098
transform 1 0 1008 0 1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_29
timestamp 1681685098
transform -1 0 1064 0 1 1370
box -8 -3 34 105
use FILL  FILL_572
timestamp 1681685098
transform 1 0 1064 0 1 1370
box -8 -3 16 105
use FILL  FILL_575
timestamp 1681685098
transform 1 0 1072 0 1 1370
box -8 -3 16 105
use FILL  FILL_577
timestamp 1681685098
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_579
timestamp 1681685098
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use FILL  FILL_581
timestamp 1681685098
transform 1 0 1096 0 1 1370
box -8 -3 16 105
use FILL  FILL_583
timestamp 1681685098
transform 1 0 1104 0 1 1370
box -8 -3 16 105
use FILL  FILL_585
timestamp 1681685098
transform 1 0 1112 0 1 1370
box -8 -3 16 105
use FILL  FILL_586
timestamp 1681685098
transform 1 0 1120 0 1 1370
box -8 -3 16 105
use FILL  FILL_587
timestamp 1681685098
transform 1 0 1128 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_30
timestamp 1681685098
transform 1 0 1136 0 1 1370
box -8 -3 34 105
use FILL  FILL_588
timestamp 1681685098
transform 1 0 1168 0 1 1370
box -8 -3 16 105
use FILL  FILL_589
timestamp 1681685098
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_590
timestamp 1681685098
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_591
timestamp 1681685098
transform 1 0 1192 0 1 1370
box -8 -3 16 105
use FILL  FILL_592
timestamp 1681685098
transform 1 0 1200 0 1 1370
box -8 -3 16 105
use FILL  FILL_593
timestamp 1681685098
transform 1 0 1208 0 1 1370
box -8 -3 16 105
use FILL  FILL_594
timestamp 1681685098
transform 1 0 1216 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_31
timestamp 1681685098
transform -1 0 1256 0 1 1370
box -8 -3 34 105
use FILL  FILL_595
timestamp 1681685098
transform 1 0 1256 0 1 1370
box -8 -3 16 105
use FILL  FILL_596
timestamp 1681685098
transform 1 0 1264 0 1 1370
box -8 -3 16 105
use FILL  FILL_597
timestamp 1681685098
transform 1 0 1272 0 1 1370
box -8 -3 16 105
use FILL  FILL_598
timestamp 1681685098
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use FILL  FILL_599
timestamp 1681685098
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_602
timestamp 1681685098
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_604
timestamp 1681685098
transform 1 0 1304 0 1 1370
box -8 -3 16 105
use FILL  FILL_605
timestamp 1681685098
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_606
timestamp 1681685098
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_28
timestamp 1681685098
transform -1 0 1352 0 1 1370
box -8 -3 32 105
use FILL  FILL_607
timestamp 1681685098
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use FILL  FILL_608
timestamp 1681685098
transform 1 0 1360 0 1 1370
box -8 -3 16 105
use FILL  FILL_609
timestamp 1681685098
transform 1 0 1368 0 1 1370
box -8 -3 16 105
use FILL  FILL_610
timestamp 1681685098
transform 1 0 1376 0 1 1370
box -8 -3 16 105
use FILL  FILL_611
timestamp 1681685098
transform 1 0 1384 0 1 1370
box -8 -3 16 105
use FILL  FILL_612
timestamp 1681685098
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_613
timestamp 1681685098
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_32
timestamp 1681685098
transform -1 0 1440 0 1 1370
box -8 -3 34 105
use FILL  FILL_614
timestamp 1681685098
transform 1 0 1440 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_10
timestamp 1681685098
transform -1 0 1480 0 1 1370
box -8 -3 40 105
use FILL  FILL_615
timestamp 1681685098
transform 1 0 1480 0 1 1370
box -8 -3 16 105
use FILL  FILL_616
timestamp 1681685098
transform 1 0 1488 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1681685098
transform -1 0 1592 0 1 1370
box -8 -3 104 105
use FILL  FILL_617
timestamp 1681685098
transform 1 0 1592 0 1 1370
box -8 -3 16 105
use FILL  FILL_623
timestamp 1681685098
transform 1 0 1600 0 1 1370
box -8 -3 16 105
use FILL  FILL_625
timestamp 1681685098
transform 1 0 1608 0 1 1370
box -8 -3 16 105
use FILL  FILL_627
timestamp 1681685098
transform 1 0 1616 0 1 1370
box -8 -3 16 105
use FILL  FILL_629
timestamp 1681685098
transform 1 0 1624 0 1 1370
box -8 -3 16 105
use FILL  FILL_631
timestamp 1681685098
transform 1 0 1632 0 1 1370
box -8 -3 16 105
use FILL  FILL_632
timestamp 1681685098
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use FILL  FILL_633
timestamp 1681685098
transform 1 0 1648 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_31
timestamp 1681685098
transform 1 0 1656 0 1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_35
timestamp 1681685098
transform 1 0 1672 0 1 1370
box -8 -3 34 105
use FILL  FILL_634
timestamp 1681685098
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_635
timestamp 1681685098
transform 1 0 1712 0 1 1370
box -8 -3 16 105
use FILL  FILL_637
timestamp 1681685098
transform 1 0 1720 0 1 1370
box -8 -3 16 105
use FILL  FILL_639
timestamp 1681685098
transform 1 0 1728 0 1 1370
box -8 -3 16 105
use FILL  FILL_640
timestamp 1681685098
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_641
timestamp 1681685098
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_642
timestamp 1681685098
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_643
timestamp 1681685098
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_644
timestamp 1681685098
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_645
timestamp 1681685098
transform 1 0 1776 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_11
timestamp 1681685098
transform 1 0 1784 0 1 1370
box -8 -3 40 105
use OR2X1  OR2X1_26
timestamp 1681685098
transform -1 0 1848 0 1 1370
box -8 -3 40 105
use FILL  FILL_646
timestamp 1681685098
transform 1 0 1848 0 1 1370
box -8 -3 16 105
use FILL  FILL_647
timestamp 1681685098
transform 1 0 1856 0 1 1370
box -8 -3 16 105
use FILL  FILL_648
timestamp 1681685098
transform 1 0 1864 0 1 1370
box -8 -3 16 105
use FILL  FILL_649
timestamp 1681685098
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use FILL  FILL_650
timestamp 1681685098
transform 1 0 1880 0 1 1370
box -8 -3 16 105
use FILL  FILL_651
timestamp 1681685098
transform 1 0 1888 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1681685098
transform -1 0 1920 0 1 1370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1681685098
transform 1 0 1920 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_32
timestamp 1681685098
transform 1 0 2016 0 1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_36
timestamp 1681685098
transform 1 0 2032 0 1 1370
box -8 -3 34 105
use FILL  FILL_652
timestamp 1681685098
transform 1 0 2064 0 1 1370
box -8 -3 16 105
use FILL  FILL_653
timestamp 1681685098
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_659
timestamp 1681685098
transform 1 0 2080 0 1 1370
box -8 -3 16 105
use FILL  FILL_661
timestamp 1681685098
transform 1 0 2088 0 1 1370
box -8 -3 16 105
use FILL  FILL_663
timestamp 1681685098
transform 1 0 2096 0 1 1370
box -8 -3 16 105
use FILL  FILL_665
timestamp 1681685098
transform 1 0 2104 0 1 1370
box -8 -3 16 105
use FILL  FILL_667
timestamp 1681685098
transform 1 0 2112 0 1 1370
box -8 -3 16 105
use FILL  FILL_669
timestamp 1681685098
transform 1 0 2120 0 1 1370
box -8 -3 16 105
use FILL  FILL_671
timestamp 1681685098
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_673
timestamp 1681685098
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_13
timestamp 1681685098
transform 1 0 2170 0 1 1370
box -10 -3 10 3
use M2_M1  M2_M1_523
timestamp 1681685098
transform 1 0 188 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1681685098
transform 1 0 84 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_386
timestamp 1681685098
transform 1 0 164 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_531
timestamp 1681685098
transform 1 0 172 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_387
timestamp 1681685098
transform 1 0 188 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_532
timestamp 1681685098
transform 1 0 196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1681685098
transform 1 0 220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1681685098
transform 1 0 116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1681685098
transform 1 0 164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1681685098
transform 1 0 180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1681685098
transform 1 0 212 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_410
timestamp 1681685098
transform 1 0 180 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_577
timestamp 1681685098
transform 1 0 236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1681685098
transform 1 0 244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1681685098
transform 1 0 220 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_411
timestamp 1681685098
transform 1 0 236 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_534
timestamp 1681685098
transform 1 0 268 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_388
timestamp 1681685098
transform 1 0 276 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_579
timestamp 1681685098
transform 1 0 276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1681685098
transform 1 0 316 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1681685098
transform 1 0 324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1681685098
transform 1 0 340 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_412
timestamp 1681685098
transform 1 0 340 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_627
timestamp 1681685098
transform 1 0 348 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_437
timestamp 1681685098
transform 1 0 340 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_537
timestamp 1681685098
transform 1 0 404 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_393
timestamp 1681685098
transform 1 0 372 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_580
timestamp 1681685098
transform 1 0 380 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_394
timestamp 1681685098
transform 1 0 396 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1681685098
transform 1 0 428 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1681685098
transform 1 0 492 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_538
timestamp 1681685098
transform 1 0 428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1681685098
transform 1 0 444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1681685098
transform 1 0 532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1681685098
transform 1 0 420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1681685098
transform 1 0 372 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1681685098
transform 1 0 396 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1681685098
transform 1 0 404 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_423
timestamp 1681685098
transform 1 0 372 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1681685098
transform 1 0 420 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_582
timestamp 1681685098
transform 1 0 492 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_374
timestamp 1681685098
transform 1 0 548 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_541
timestamp 1681685098
transform 1 0 548 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_360
timestamp 1681685098
transform 1 0 572 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_542
timestamp 1681685098
transform 1 0 572 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1681685098
transform 1 0 548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1681685098
transform 1 0 564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1681685098
transform 1 0 548 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_395
timestamp 1681685098
transform 1 0 588 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1681685098
transform 1 0 580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1681685098
transform 1 0 572 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_585
timestamp 1681685098
transform 1 0 628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1681685098
transform 1 0 612 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_414
timestamp 1681685098
transform 1 0 620 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_628
timestamp 1681685098
transform 1 0 620 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1681685098
transform 1 0 644 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_425
timestamp 1681685098
transform 1 0 644 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_586
timestamp 1681685098
transform 1 0 660 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_375
timestamp 1681685098
transform 1 0 692 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_525
timestamp 1681685098
transform 1 0 700 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1681685098
transform 1 0 692 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_445
timestamp 1681685098
transform 1 0 676 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_587
timestamp 1681685098
transform 1 0 708 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_426
timestamp 1681685098
transform 1 0 708 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_544
timestamp 1681685098
transform 1 0 740 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_367
timestamp 1681685098
transform 1 0 804 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1681685098
transform 1 0 780 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_545
timestamp 1681685098
transform 1 0 756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1681685098
transform 1 0 780 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_415
timestamp 1681685098
transform 1 0 756 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_547
timestamp 1681685098
transform 1 0 828 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_396
timestamp 1681685098
transform 1 0 804 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1681685098
transform 1 0 796 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_588
timestamp 1681685098
transform 1 0 836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1681685098
transform 1 0 836 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1681685098
transform 1 0 892 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_397
timestamp 1681685098
transform 1 0 900 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1681685098
transform 1 0 892 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_629
timestamp 1681685098
transform 1 0 900 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1681685098
transform 1 0 916 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1681685098
transform 1 0 916 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_377
timestamp 1681685098
transform 1 0 948 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1681685098
transform 1 0 964 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_549
timestamp 1681685098
transform 1 0 956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1681685098
transform 1 0 948 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_398
timestamp 1681685098
transform 1 0 956 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_619
timestamp 1681685098
transform 1 0 956 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1681685098
transform 1 0 1020 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1681685098
transform 1 0 1044 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_427
timestamp 1681685098
transform 1 0 1028 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_550
timestamp 1681685098
transform 1 0 1060 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_399
timestamp 1681685098
transform 1 0 1052 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1681685098
transform 1 0 1068 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_621
timestamp 1681685098
transform 1 0 1076 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1681685098
transform 1 0 1068 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_438
timestamp 1681685098
transform 1 0 1068 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1681685098
transform 1 0 1100 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1681685098
transform 1 0 1116 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1681685098
transform 1 0 1212 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1681685098
transform 1 0 1140 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1681685098
transform 1 0 1132 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1681685098
transform 1 0 1228 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_527
timestamp 1681685098
transform 1 0 1244 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_390
timestamp 1681685098
transform 1 0 1164 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_551
timestamp 1681685098
transform 1 0 1228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1681685098
transform 1 0 1132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1681685098
transform 1 0 1148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1681685098
transform 1 0 1180 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_428
timestamp 1681685098
transform 1 0 1156 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1681685098
transform 1 0 1140 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1681685098
transform 1 0 1148 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_552
timestamp 1681685098
transform 1 0 1252 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1681685098
transform 1 0 1260 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_401
timestamp 1681685098
transform 1 0 1252 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_594
timestamp 1681685098
transform 1 0 1260 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_402
timestamp 1681685098
transform 1 0 1268 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_595
timestamp 1681685098
transform 1 0 1276 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_440
timestamp 1681685098
transform 1 0 1260 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1681685098
transform 1 0 1292 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_554
timestamp 1681685098
transform 1 0 1292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1681685098
transform 1 0 1284 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_429
timestamp 1681685098
transform 1 0 1284 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_555
timestamp 1681685098
transform 1 0 1364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1681685098
transform 1 0 1372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1681685098
transform 1 0 1332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1681685098
transform 1 0 1340 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_403
timestamp 1681685098
transform 1 0 1364 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1681685098
transform 1 0 1468 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1681685098
transform 1 0 1452 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1681685098
transform 1 0 1412 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_557
timestamp 1681685098
transform 1 0 1396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1681685098
transform 1 0 1412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1681685098
transform 1 0 1380 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_404
timestamp 1681685098
transform 1 0 1396 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1681685098
transform 1 0 1500 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_559
timestamp 1681685098
transform 1 0 1508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1681685098
transform 1 0 1436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1681685098
transform 1 0 1492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1681685098
transform 1 0 1500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1681685098
transform 1 0 1396 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_430
timestamp 1681685098
transform 1 0 1380 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1681685098
transform 1 0 1492 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1681685098
transform 1 0 1508 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1681685098
transform 1 0 1500 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1681685098
transform 1 0 1540 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_560
timestamp 1681685098
transform 1 0 1540 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_381
timestamp 1681685098
transform 1 0 1580 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_561
timestamp 1681685098
transform 1 0 1564 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1681685098
transform 1 0 1548 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_405
timestamp 1681685098
transform 1 0 1556 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_624
timestamp 1681685098
transform 1 0 1572 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_432
timestamp 1681685098
transform 1 0 1572 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_562
timestamp 1681685098
transform 1 0 1604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1681685098
transform 1 0 1612 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_406
timestamp 1681685098
transform 1 0 1612 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1681685098
transform 1 0 1676 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_564
timestamp 1681685098
transform 1 0 1684 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1681685098
transform 1 0 1708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1681685098
transform 1 0 1700 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_407
timestamp 1681685098
transform 1 0 1708 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_625
timestamp 1681685098
transform 1 0 1724 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_433
timestamp 1681685098
transform 1 0 1724 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1681685098
transform 1 0 1780 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_528
timestamp 1681685098
transform 1 0 1788 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_372
timestamp 1681685098
transform 1 0 1804 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_566
timestamp 1681685098
transform 1 0 1780 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1681685098
transform 1 0 1788 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1681685098
transform 1 0 1764 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_391
timestamp 1681685098
transform 1 0 1796 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1681685098
transform 1 0 1788 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1681685098
transform 1 0 1780 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1681685098
transform 1 0 1756 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1681685098
transform 1 0 1836 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1681685098
transform 1 0 1828 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_568
timestamp 1681685098
transform 1 0 1836 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1681685098
transform 1 0 1820 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1681685098
transform 1 0 1828 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_421
timestamp 1681685098
transform 1 0 1844 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_569
timestamp 1681685098
transform 1 0 1932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1681685098
transform 1 0 1884 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_422
timestamp 1681685098
transform 1 0 1884 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1681685098
transform 1 0 1908 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1681685098
transform 1 0 1940 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1681685098
transform 1 0 1964 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_570
timestamp 1681685098
transform 1 0 1964 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_365
timestamp 1681685098
transform 1 0 2012 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_571
timestamp 1681685098
transform 1 0 2012 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_409
timestamp 1681685098
transform 1 0 1988 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1681685098
transform 1 0 2044 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1681685098
transform 1 0 2036 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_529
timestamp 1681685098
transform 1 0 2044 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1681685098
transform 1 0 2036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1681685098
transform 1 0 2028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1681685098
transform 1 0 2036 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_442
timestamp 1681685098
transform 1 0 2036 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1681685098
transform 1 0 2060 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_609
timestamp 1681685098
transform 1 0 2140 0 1 1325
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_14
timestamp 1681685098
transform 1 0 24 0 1 1270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_25
timestamp 1681685098
transform 1 0 72 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_24
timestamp 1681685098
transform 1 0 168 0 -1 1370
box -9 -3 26 105
use OR2X1  OR2X1_23
timestamp 1681685098
transform 1 0 184 0 -1 1370
box -8 -3 40 105
use OAI21X1  OAI21X1_25
timestamp 1681685098
transform -1 0 248 0 -1 1370
box -8 -3 34 105
use FILL  FILL_497
timestamp 1681685098
transform 1 0 248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_499
timestamp 1681685098
transform 1 0 256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_501
timestamp 1681685098
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_505
timestamp 1681685098
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_7
timestamp 1681685098
transform -1 0 304 0 -1 1370
box -8 -3 32 105
use FILL  FILL_506
timestamp 1681685098
transform 1 0 304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_508
timestamp 1681685098
transform 1 0 312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_522
timestamp 1681685098
transform 1 0 320 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_26
timestamp 1681685098
transform -1 0 344 0 -1 1370
box -9 -3 26 105
use FILL  FILL_523
timestamp 1681685098
transform 1 0 344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_524
timestamp 1681685098
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_525
timestamp 1681685098
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_7
timestamp 1681685098
transform 1 0 368 0 -1 1370
box -8 -3 40 105
use OAI21X1  OAI21X1_26
timestamp 1681685098
transform -1 0 432 0 -1 1370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1681685098
transform 1 0 432 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_27
timestamp 1681685098
transform 1 0 528 0 -1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_27
timestamp 1681685098
transform -1 0 576 0 -1 1370
box -8 -3 34 105
use FILL  FILL_526
timestamp 1681685098
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_528
timestamp 1681685098
transform 1 0 584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_530
timestamp 1681685098
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_537
timestamp 1681685098
transform 1 0 600 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_8
timestamp 1681685098
transform -1 0 640 0 -1 1370
box -8 -3 40 105
use FILL  FILL_538
timestamp 1681685098
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_540
timestamp 1681685098
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_542
timestamp 1681685098
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_549
timestamp 1681685098
transform 1 0 664 0 -1 1370
box -8 -3 16 105
use OR2X1  OR2X1_24
timestamp 1681685098
transform -1 0 704 0 -1 1370
box -8 -3 40 105
use INVX2  INVX2_29
timestamp 1681685098
transform -1 0 720 0 -1 1370
box -9 -3 26 105
use FILL  FILL_550
timestamp 1681685098
transform 1 0 720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_551
timestamp 1681685098
transform 1 0 728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_552
timestamp 1681685098
transform 1 0 736 0 -1 1370
box -8 -3 16 105
use OR2X1  OR2X1_25
timestamp 1681685098
transform 1 0 744 0 -1 1370
box -8 -3 40 105
use XNOR2X1  XNOR2X1_24
timestamp 1681685098
transform 1 0 776 0 -1 1370
box -8 -3 64 105
use FILL  FILL_553
timestamp 1681685098
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_554
timestamp 1681685098
transform 1 0 840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_556
timestamp 1681685098
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_557
timestamp 1681685098
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_558
timestamp 1681685098
transform 1 0 864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_559
timestamp 1681685098
transform 1 0 872 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_9
timestamp 1681685098
transform 1 0 880 0 -1 1370
box -8 -3 40 105
use FILL  FILL_560
timestamp 1681685098
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_561
timestamp 1681685098
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_562
timestamp 1681685098
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_23
timestamp 1681685098
transform 1 0 936 0 -1 1370
box -8 -3 32 105
use FILL  FILL_563
timestamp 1681685098
transform 1 0 960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_564
timestamp 1681685098
transform 1 0 968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_565
timestamp 1681685098
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_567
timestamp 1681685098
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_569
timestamp 1681685098
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_571
timestamp 1681685098
transform 1 0 1000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_573
timestamp 1681685098
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_25
timestamp 1681685098
transform -1 0 1040 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1681685098
transform 1 0 1040 0 -1 1370
box -8 -3 32 105
use FILL  FILL_574
timestamp 1681685098
transform 1 0 1064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_576
timestamp 1681685098
transform 1 0 1072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_578
timestamp 1681685098
transform 1 0 1080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_580
timestamp 1681685098
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_582
timestamp 1681685098
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_584
timestamp 1681685098
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_600
timestamp 1681685098
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_26
timestamp 1681685098
transform -1 0 1144 0 -1 1370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1681685098
transform -1 0 1240 0 -1 1370
box -8 -3 104 105
use NOR2X1  NOR2X1_9
timestamp 1681685098
transform 1 0 1240 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1681685098
transform 1 0 1264 0 -1 1370
box -8 -3 32 105
use FILL  FILL_601
timestamp 1681685098
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_603
timestamp 1681685098
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_618
timestamp 1681685098
transform 1 0 1304 0 -1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_0
timestamp 1681685098
transform -1 0 1368 0 -1 1370
box -8 -3 64 105
use OAI21X1  OAI21X1_33
timestamp 1681685098
transform 1 0 1368 0 -1 1370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1681685098
transform 1 0 1400 0 -1 1370
box -8 -3 104 105
use FILL  FILL_619
timestamp 1681685098
transform 1 0 1496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_620
timestamp 1681685098
transform 1 0 1504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_621
timestamp 1681685098
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_30
timestamp 1681685098
transform 1 0 1520 0 -1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_34
timestamp 1681685098
transform 1 0 1536 0 -1 1370
box -8 -3 34 105
use NAND2X1  NAND2X1_29
timestamp 1681685098
transform -1 0 1592 0 -1 1370
box -8 -3 32 105
use M3_M2  M3_M2_448
timestamp 1681685098
transform 1 0 1604 0 1 1275
box -3 -3 3 3
use FILL  FILL_622
timestamp 1681685098
transform 1 0 1592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_624
timestamp 1681685098
transform 1 0 1600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_626
timestamp 1681685098
transform 1 0 1608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_628
timestamp 1681685098
transform 1 0 1616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_630
timestamp 1681685098
transform 1 0 1624 0 -1 1370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_25
timestamp 1681685098
transform 1 0 1632 0 -1 1370
box -8 -3 64 105
use NAND2X1  NAND2X1_30
timestamp 1681685098
transform 1 0 1688 0 -1 1370
box -8 -3 32 105
use FILL  FILL_636
timestamp 1681685098
transform 1 0 1712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_638
timestamp 1681685098
transform 1 0 1720 0 -1 1370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_26
timestamp 1681685098
transform 1 0 1728 0 -1 1370
box -8 -3 64 105
use FILL  FILL_654
timestamp 1681685098
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use OR2X1  OR2X1_27
timestamp 1681685098
transform 1 0 1792 0 -1 1370
box -8 -3 40 105
use INVX2  INVX2_33
timestamp 1681685098
transform -1 0 1840 0 -1 1370
box -9 -3 26 105
use FILL  FILL_655
timestamp 1681685098
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1681685098
transform -1 0 1944 0 -1 1370
box -8 -3 104 105
use FILL  FILL_656
timestamp 1681685098
transform 1 0 1944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_657
timestamp 1681685098
transform 1 0 1952 0 -1 1370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_27
timestamp 1681685098
transform 1 0 1960 0 -1 1370
box -8 -3 64 105
use NAND2X1  NAND2X1_31
timestamp 1681685098
transform 1 0 2016 0 -1 1370
box -8 -3 32 105
use OR2X1  OR2X1_28
timestamp 1681685098
transform 1 0 2040 0 -1 1370
box -8 -3 40 105
use FILL  FILL_658
timestamp 1681685098
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_660
timestamp 1681685098
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_662
timestamp 1681685098
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_664
timestamp 1681685098
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_666
timestamp 1681685098
transform 1 0 2104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_668
timestamp 1681685098
transform 1 0 2112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_670
timestamp 1681685098
transform 1 0 2120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_672
timestamp 1681685098
transform 1 0 2128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_674
timestamp 1681685098
transform 1 0 2136 0 -1 1370
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_15
timestamp 1681685098
transform 1 0 2194 0 1 1270
box -10 -3 10 3
use M3_M2  M3_M2_451
timestamp 1681685098
transform 1 0 92 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_637
timestamp 1681685098
transform 1 0 100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1681685098
transform 1 0 148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1681685098
transform 1 0 156 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_456
timestamp 1681685098
transform 1 0 212 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_631
timestamp 1681685098
transform 1 0 212 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_452
timestamp 1681685098
transform 1 0 244 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1681685098
transform 1 0 260 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1681685098
transform 1 0 252 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1681685098
transform 1 0 228 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_681
timestamp 1681685098
transform 1 0 204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1681685098
transform 1 0 228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1681685098
transform 1 0 236 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_461
timestamp 1681685098
transform 1 0 268 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1681685098
transform 1 0 316 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_639
timestamp 1681685098
transform 1 0 268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1681685098
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_466
timestamp 1681685098
transform 1 0 292 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_641
timestamp 1681685098
transform 1 0 316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1681685098
transform 1 0 340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1681685098
transform 1 0 396 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1681685098
transform 1 0 260 0 1 1207
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1681685098
transform 1 0 268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1681685098
transform 1 0 316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1681685098
transform 1 0 324 0 1 1207
box -2 -2 2 2
use M3_M2  M3_M2_467
timestamp 1681685098
transform 1 0 420 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_686
timestamp 1681685098
transform 1 0 420 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_468
timestamp 1681685098
transform 1 0 444 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_644
timestamp 1681685098
transform 1 0 476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1681685098
transform 1 0 532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1681685098
transform 1 0 564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1681685098
transform 1 0 588 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_449
timestamp 1681685098
transform 1 0 628 0 1 1265
box -3 -3 3 3
use M2_M1  M2_M1_688
timestamp 1681685098
transform 1 0 612 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1681685098
transform 1 0 636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1681685098
transform 1 0 644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1681685098
transform 1 0 676 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_480
timestamp 1681685098
transform 1 0 676 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_690
timestamp 1681685098
transform 1 0 708 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_458
timestamp 1681685098
transform 1 0 732 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_632
timestamp 1681685098
transform 1 0 732 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_459
timestamp 1681685098
transform 1 0 788 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1681685098
transform 1 0 756 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_648
timestamp 1681685098
transform 1 0 756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1681685098
transform 1 0 788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1681685098
transform 1 0 740 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1681685098
transform 1 0 796 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_464
timestamp 1681685098
transform 1 0 820 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_650
timestamp 1681685098
transform 1 0 820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1681685098
transform 1 0 796 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_481
timestamp 1681685098
transform 1 0 812 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1681685098
transform 1 0 796 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1681685098
transform 1 0 836 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1681685098
transform 1 0 844 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_693
timestamp 1681685098
transform 1 0 860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1681685098
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1681685098
transform 1 0 916 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_482
timestamp 1681685098
transform 1 0 924 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_652
timestamp 1681685098
transform 1 0 948 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1681685098
transform 1 0 964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1681685098
transform 1 0 964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1681685098
transform 1 0 1020 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1681685098
transform 1 0 1028 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1681685098
transform 1 0 1068 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1681685098
transform 1 0 1052 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1681685098
transform 1 0 1060 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1681685098
transform 1 0 1084 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_474
timestamp 1681685098
transform 1 0 1108 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_655
timestamp 1681685098
transform 1 0 1148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1681685098
transform 1 0 1140 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_475
timestamp 1681685098
transform 1 0 1148 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_656
timestamp 1681685098
transform 1 0 1180 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1681685098
transform 1 0 1188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1681685098
transform 1 0 1196 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1681685098
transform 1 0 1172 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_483
timestamp 1681685098
transform 1 0 1140 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1681685098
transform 1 0 1180 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1681685098
transform 1 0 1196 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_715
timestamp 1681685098
transform 1 0 1284 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_454
timestamp 1681685098
transform 1 0 1316 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1681685098
transform 1 0 1340 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1681685098
transform 1 0 1332 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_659
timestamp 1681685098
transform 1 0 1340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1681685098
transform 1 0 1356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1681685098
transform 1 0 1364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1681685098
transform 1 0 1324 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1681685098
transform 1 0 1332 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_470
timestamp 1681685098
transform 1 0 1372 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_662
timestamp 1681685098
transform 1 0 1380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1681685098
transform 1 0 1396 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1681685098
transform 1 0 1452 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_486
timestamp 1681685098
transform 1 0 1452 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_664
timestamp 1681685098
transform 1 0 1468 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1681685098
transform 1 0 1564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1681685098
transform 1 0 1604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1681685098
transform 1 0 1524 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_487
timestamp 1681685098
transform 1 0 1524 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_705
timestamp 1681685098
transform 1 0 1612 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_476
timestamp 1681685098
transform 1 0 1652 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_716
timestamp 1681685098
transform 1 0 1652 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_477
timestamp 1681685098
transform 1 0 1684 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_667
timestamp 1681685098
transform 1 0 1708 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1681685098
transform 1 0 1724 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1681685098
transform 1 0 1764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1681685098
transform 1 0 1748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1681685098
transform 1 0 1756 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_478
timestamp 1681685098
transform 1 0 1764 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_635
timestamp 1681685098
transform 1 0 1780 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_460
timestamp 1681685098
transform 1 0 1828 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_636
timestamp 1681685098
transform 1 0 1836 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1681685098
transform 1 0 1812 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1681685098
transform 1 0 1820 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_471
timestamp 1681685098
transform 1 0 1828 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_708
timestamp 1681685098
transform 1 0 1804 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_479
timestamp 1681685098
transform 1 0 1812 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_672
timestamp 1681685098
transform 1 0 1844 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_472
timestamp 1681685098
transform 1 0 1860 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_673
timestamp 1681685098
transform 1 0 1884 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_473
timestamp 1681685098
transform 1 0 1932 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_674
timestamp 1681685098
transform 1 0 1940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1681685098
transform 1 0 1860 0 1 1207
box -2 -2 2 2
use M3_M2  M3_M2_488
timestamp 1681685098
transform 1 0 1940 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_709
timestamp 1681685098
transform 1 0 1956 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1681685098
transform 1 0 1948 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_492
timestamp 1681685098
transform 1 0 1948 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_675
timestamp 1681685098
transform 1 0 1988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1681685098
transform 1 0 1972 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1681685098
transform 1 0 1996 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1681685098
transform 1 0 2052 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1681685098
transform 1 0 2044 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_489
timestamp 1681685098
transform 1 0 2044 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1681685098
transform 1 0 2012 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1681685098
transform 1 0 2028 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1681685098
transform 1 0 2052 0 1 1185
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_16
timestamp 1681685098
transform 1 0 48 0 1 1170
box -10 -3 10 3
use FILL  FILL_675
timestamp 1681685098
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_677
timestamp 1681685098
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_679
timestamp 1681685098
transform 1 0 88 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_34
timestamp 1681685098
transform -1 0 112 0 1 1170
box -9 -3 26 105
use FILL  FILL_680
timestamp 1681685098
transform 1 0 112 0 1 1170
box -8 -3 16 105
use FILL  FILL_681
timestamp 1681685098
transform 1 0 120 0 1 1170
box -8 -3 16 105
use FILL  FILL_683
timestamp 1681685098
transform 1 0 128 0 1 1170
box -8 -3 16 105
use FILL  FILL_685
timestamp 1681685098
transform 1 0 136 0 1 1170
box -8 -3 16 105
use FILL  FILL_686
timestamp 1681685098
transform 1 0 144 0 1 1170
box -8 -3 16 105
use XNOR2X1  XNOR2X1_28
timestamp 1681685098
transform -1 0 208 0 1 1170
box -8 -3 64 105
use NAND2X1  NAND2X1_32
timestamp 1681685098
transform -1 0 232 0 1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_38
timestamp 1681685098
transform -1 0 264 0 1 1170
box -8 -3 34 105
use XNOR2X1  XNOR2X1_29
timestamp 1681685098
transform -1 0 320 0 1 1170
box -8 -3 64 105
use INVX2  INVX2_35
timestamp 1681685098
transform 1 0 320 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1681685098
transform -1 0 432 0 1 1170
box -8 -3 104 105
use FILL  FILL_687
timestamp 1681685098
transform 1 0 432 0 1 1170
box -8 -3 16 105
use FILL  FILL_688
timestamp 1681685098
transform 1 0 440 0 1 1170
box -8 -3 16 105
use FILL  FILL_689
timestamp 1681685098
transform 1 0 448 0 1 1170
box -8 -3 16 105
use FILL  FILL_690
timestamp 1681685098
transform 1 0 456 0 1 1170
box -8 -3 16 105
use FILL  FILL_691
timestamp 1681685098
transform 1 0 464 0 1 1170
box -8 -3 16 105
use FILL  FILL_692
timestamp 1681685098
transform 1 0 472 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1681685098
transform -1 0 576 0 1 1170
box -8 -3 104 105
use FILL  FILL_693
timestamp 1681685098
transform 1 0 576 0 1 1170
box -8 -3 16 105
use FILL  FILL_703
timestamp 1681685098
transform 1 0 584 0 1 1170
box -8 -3 16 105
use FILL  FILL_705
timestamp 1681685098
transform 1 0 592 0 1 1170
box -8 -3 16 105
use FILL  FILL_707
timestamp 1681685098
transform 1 0 600 0 1 1170
box -8 -3 16 105
use OR2X1  OR2X1_29
timestamp 1681685098
transform 1 0 608 0 1 1170
box -8 -3 40 105
use FILL  FILL_708
timestamp 1681685098
transform 1 0 640 0 1 1170
box -8 -3 16 105
use FILL  FILL_711
timestamp 1681685098
transform 1 0 648 0 1 1170
box -8 -3 16 105
use FILL  FILL_713
timestamp 1681685098
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_715
timestamp 1681685098
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_716
timestamp 1681685098
transform 1 0 672 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_40
timestamp 1681685098
transform 1 0 680 0 1 1170
box -8 -3 34 105
use FILL  FILL_717
timestamp 1681685098
transform 1 0 712 0 1 1170
box -8 -3 16 105
use FILL  FILL_718
timestamp 1681685098
transform 1 0 720 0 1 1170
box -8 -3 16 105
use FILL  FILL_719
timestamp 1681685098
transform 1 0 728 0 1 1170
box -8 -3 16 105
use XNOR2X1  XNOR2X1_30
timestamp 1681685098
transform -1 0 792 0 1 1170
box -8 -3 64 105
use AOI21X1  AOI21X1_3
timestamp 1681685098
transform -1 0 824 0 1 1170
box -7 -3 39 105
use FILL  FILL_720
timestamp 1681685098
transform 1 0 824 0 1 1170
box -8 -3 16 105
use FILL  FILL_724
timestamp 1681685098
transform 1 0 832 0 1 1170
box -8 -3 16 105
use FILL  FILL_726
timestamp 1681685098
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_727
timestamp 1681685098
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_728
timestamp 1681685098
transform 1 0 856 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_38
timestamp 1681685098
transform 1 0 864 0 1 1170
box -9 -3 26 105
use FILL  FILL_729
timestamp 1681685098
transform 1 0 880 0 1 1170
box -8 -3 16 105
use FILL  FILL_730
timestamp 1681685098
transform 1 0 888 0 1 1170
box -8 -3 16 105
use FILL  FILL_732
timestamp 1681685098
transform 1 0 896 0 1 1170
box -8 -3 16 105
use FILL  FILL_734
timestamp 1681685098
transform 1 0 904 0 1 1170
box -8 -3 16 105
use FILL  FILL_736
timestamp 1681685098
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_738
timestamp 1681685098
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_740
timestamp 1681685098
transform 1 0 928 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_41
timestamp 1681685098
transform 1 0 936 0 1 1170
box -8 -3 34 105
use FILL  FILL_742
timestamp 1681685098
transform 1 0 968 0 1 1170
box -8 -3 16 105
use FILL  FILL_748
timestamp 1681685098
transform 1 0 976 0 1 1170
box -8 -3 16 105
use FILL  FILL_750
timestamp 1681685098
transform 1 0 984 0 1 1170
box -8 -3 16 105
use FILL  FILL_752
timestamp 1681685098
transform 1 0 992 0 1 1170
box -8 -3 16 105
use FILL  FILL_754
timestamp 1681685098
transform 1 0 1000 0 1 1170
box -8 -3 16 105
use FILL  FILL_756
timestamp 1681685098
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use FILL  FILL_757
timestamp 1681685098
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_34
timestamp 1681685098
transform -1 0 1048 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1681685098
transform 1 0 1048 0 1 1170
box -8 -3 32 105
use FILL  FILL_758
timestamp 1681685098
transform 1 0 1072 0 1 1170
box -8 -3 16 105
use FILL  FILL_762
timestamp 1681685098
transform 1 0 1080 0 1 1170
box -8 -3 16 105
use FILL  FILL_764
timestamp 1681685098
transform 1 0 1088 0 1 1170
box -8 -3 16 105
use FILL  FILL_766
timestamp 1681685098
transform 1 0 1096 0 1 1170
box -8 -3 16 105
use FILL  FILL_768
timestamp 1681685098
transform 1 0 1104 0 1 1170
box -8 -3 16 105
use FILL  FILL_769
timestamp 1681685098
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_770
timestamp 1681685098
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use FILL  FILL_771
timestamp 1681685098
transform 1 0 1128 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_496
timestamp 1681685098
transform 1 0 1172 0 1 1175
box -3 -3 3 3
use AND2X2  AND2X2_1
timestamp 1681685098
transform 1 0 1136 0 1 1170
box -8 -3 40 105
use FILL  FILL_772
timestamp 1681685098
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_497
timestamp 1681685098
transform 1 0 1228 0 1 1175
box -3 -3 3 3
use FAX1  FAX1_0
timestamp 1681685098
transform 1 0 1176 0 1 1170
box -5 -3 126 105
use FILL  FILL_775
timestamp 1681685098
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_776
timestamp 1681685098
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use FILL  FILL_777
timestamp 1681685098
transform 1 0 1312 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_498
timestamp 1681685098
transform 1 0 1340 0 1 1175
box -3 -3 3 3
use FILL  FILL_778
timestamp 1681685098
transform 1 0 1320 0 1 1170
box -8 -3 16 105
use AND2X2  AND2X2_2
timestamp 1681685098
transform 1 0 1328 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1681685098
transform -1 0 1392 0 1 1170
box -8 -3 40 105
use FILL  FILL_779
timestamp 1681685098
transform 1 0 1392 0 1 1170
box -8 -3 16 105
use FILL  FILL_780
timestamp 1681685098
transform 1 0 1400 0 1 1170
box -8 -3 16 105
use FILL  FILL_781
timestamp 1681685098
transform 1 0 1408 0 1 1170
box -8 -3 16 105
use FILL  FILL_791
timestamp 1681685098
transform 1 0 1416 0 1 1170
box -8 -3 16 105
use FILL  FILL_793
timestamp 1681685098
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use FILL  FILL_795
timestamp 1681685098
transform 1 0 1432 0 1 1170
box -8 -3 16 105
use FILL  FILL_797
timestamp 1681685098
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use BUFX2  BUFX2_3
timestamp 1681685098
transform -1 0 1472 0 1 1170
box -5 -3 28 105
use FILL  FILL_798
timestamp 1681685098
transform 1 0 1472 0 1 1170
box -8 -3 16 105
use FILL  FILL_799
timestamp 1681685098
transform 1 0 1480 0 1 1170
box -8 -3 16 105
use FILL  FILL_800
timestamp 1681685098
transform 1 0 1488 0 1 1170
box -8 -3 16 105
use FILL  FILL_801
timestamp 1681685098
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use FILL  FILL_802
timestamp 1681685098
transform 1 0 1504 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1681685098
transform 1 0 1512 0 1 1170
box -8 -3 104 105
use FILL  FILL_803
timestamp 1681685098
transform 1 0 1608 0 1 1170
box -8 -3 16 105
use FILL  FILL_817
timestamp 1681685098
transform 1 0 1616 0 1 1170
box -8 -3 16 105
use FILL  FILL_819
timestamp 1681685098
transform 1 0 1624 0 1 1170
box -8 -3 16 105
use FILL  FILL_821
timestamp 1681685098
transform 1 0 1632 0 1 1170
box -8 -3 16 105
use FILL  FILL_823
timestamp 1681685098
transform 1 0 1640 0 1 1170
box -8 -3 16 105
use OR2X1  OR2X1_31
timestamp 1681685098
transform 1 0 1648 0 1 1170
box -8 -3 40 105
use FILL  FILL_824
timestamp 1681685098
transform 1 0 1680 0 1 1170
box -8 -3 16 105
use FILL  FILL_829
timestamp 1681685098
transform 1 0 1688 0 1 1170
box -8 -3 16 105
use FILL  FILL_831
timestamp 1681685098
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_833
timestamp 1681685098
transform 1 0 1704 0 1 1170
box -8 -3 16 105
use FILL  FILL_835
timestamp 1681685098
transform 1 0 1712 0 1 1170
box -8 -3 16 105
use FILL  FILL_836
timestamp 1681685098
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use OR2X1  OR2X1_32
timestamp 1681685098
transform -1 0 1760 0 1 1170
box -8 -3 40 105
use NAND2X1  NAND2X1_35
timestamp 1681685098
transform 1 0 1760 0 1 1170
box -8 -3 32 105
use FILL  FILL_837
timestamp 1681685098
transform 1 0 1784 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_499
timestamp 1681685098
transform 1 0 1804 0 1 1175
box -3 -3 3 3
use FILL  FILL_842
timestamp 1681685098
transform 1 0 1792 0 1 1170
box -8 -3 16 105
use FILL  FILL_844
timestamp 1681685098
transform 1 0 1800 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_43
timestamp 1681685098
transform 1 0 1808 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_500
timestamp 1681685098
transform 1 0 1852 0 1 1175
box -3 -3 3 3
use FILL  FILL_846
timestamp 1681685098
transform 1 0 1840 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1681685098
transform 1 0 1848 0 1 1170
box -8 -3 104 105
use FILL  FILL_847
timestamp 1681685098
transform 1 0 1944 0 1 1170
box -8 -3 16 105
use FILL  FILL_848
timestamp 1681685098
transform 1 0 1952 0 1 1170
box -8 -3 16 105
use OR2X1  OR2X1_33
timestamp 1681685098
transform 1 0 1960 0 1 1170
box -8 -3 40 105
use XNOR2X1  XNOR2X1_31
timestamp 1681685098
transform 1 0 1992 0 1 1170
box -8 -3 64 105
use FILL  FILL_849
timestamp 1681685098
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_858
timestamp 1681685098
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use FILL  FILL_860
timestamp 1681685098
transform 1 0 2064 0 1 1170
box -8 -3 16 105
use FILL  FILL_862
timestamp 1681685098
transform 1 0 2072 0 1 1170
box -8 -3 16 105
use FILL  FILL_864
timestamp 1681685098
transform 1 0 2080 0 1 1170
box -8 -3 16 105
use FILL  FILL_866
timestamp 1681685098
transform 1 0 2088 0 1 1170
box -8 -3 16 105
use FILL  FILL_868
timestamp 1681685098
transform 1 0 2096 0 1 1170
box -8 -3 16 105
use FILL  FILL_870
timestamp 1681685098
transform 1 0 2104 0 1 1170
box -8 -3 16 105
use FILL  FILL_872
timestamp 1681685098
transform 1 0 2112 0 1 1170
box -8 -3 16 105
use FILL  FILL_874
timestamp 1681685098
transform 1 0 2120 0 1 1170
box -8 -3 16 105
use FILL  FILL_876
timestamp 1681685098
transform 1 0 2128 0 1 1170
box -8 -3 16 105
use FILL  FILL_878
timestamp 1681685098
transform 1 0 2136 0 1 1170
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_17
timestamp 1681685098
transform 1 0 2170 0 1 1170
box -10 -3 10 3
use M2_M1  M2_M1_722
timestamp 1681685098
transform 1 0 84 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1681685098
transform 1 0 116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1681685098
transform 1 0 100 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_505
timestamp 1681685098
transform 1 0 140 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_802
timestamp 1681685098
transform 1 0 140 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_506
timestamp 1681685098
transform 1 0 212 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_724
timestamp 1681685098
transform 1 0 164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1681685098
transform 1 0 172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1681685098
transform 1 0 164 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_513
timestamp 1681685098
transform 1 0 236 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1681685098
transform 1 0 260 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_726
timestamp 1681685098
transform 1 0 220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1681685098
transform 1 0 236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1681685098
transform 1 0 260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1681685098
transform 1 0 316 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_528
timestamp 1681685098
transform 1 0 220 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1681685098
transform 1 0 236 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_766
timestamp 1681685098
transform 1 0 340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1681685098
transform 1 0 356 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_529
timestamp 1681685098
transform 1 0 356 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1681685098
transform 1 0 404 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_728
timestamp 1681685098
transform 1 0 404 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_507
timestamp 1681685098
transform 1 0 492 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1681685098
transform 1 0 476 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_729
timestamp 1681685098
transform 1 0 492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1681685098
transform 1 0 508 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1681685098
transform 1 0 412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1681685098
transform 1 0 468 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_530
timestamp 1681685098
transform 1 0 412 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1681685098
transform 1 0 444 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1681685098
transform 1 0 420 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_731
timestamp 1681685098
transform 1 0 532 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_517
timestamp 1681685098
transform 1 0 548 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_732
timestamp 1681685098
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1681685098
transform 1 0 516 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1681685098
transform 1 0 532 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_524
timestamp 1681685098
transform 1 0 540 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_772
timestamp 1681685098
transform 1 0 548 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1681685098
transform 1 0 532 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_508
timestamp 1681685098
transform 1 0 564 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_733
timestamp 1681685098
transform 1 0 580 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1681685098
transform 1 0 628 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_509
timestamp 1681685098
transform 1 0 660 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_734
timestamp 1681685098
transform 1 0 660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1681685098
transform 1 0 676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1681685098
transform 1 0 788 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1681685098
transform 1 0 772 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1681685098
transform 1 0 708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1681685098
transform 1 0 756 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1681685098
transform 1 0 764 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_532
timestamp 1681685098
transform 1 0 676 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1681685098
transform 1 0 748 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_777
timestamp 1681685098
transform 1 0 788 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_541
timestamp 1681685098
transform 1 0 764 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1681685098
transform 1 0 780 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1681685098
transform 1 0 804 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_737
timestamp 1681685098
transform 1 0 804 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1681685098
transform 1 0 804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1681685098
transform 1 0 812 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_534
timestamp 1681685098
transform 1 0 804 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1681685098
transform 1 0 844 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_738
timestamp 1681685098
transform 1 0 844 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_520
timestamp 1681685098
transform 1 0 876 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_719
timestamp 1681685098
transform 1 0 884 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1681685098
transform 1 0 876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1681685098
transform 1 0 860 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1681685098
transform 1 0 892 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1681685098
transform 1 0 1036 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1681685098
transform 1 0 1028 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_525
timestamp 1681685098
transform 1 0 1036 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_804
timestamp 1681685098
transform 1 0 1036 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1681685098
transform 1 0 1060 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1681685098
transform 1 0 1076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1681685098
transform 1 0 1108 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_526
timestamp 1681685098
transform 1 0 1108 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_784
timestamp 1681685098
transform 1 0 1132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_501
timestamp 1681685098
transform 1 0 1172 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_743
timestamp 1681685098
transform 1 0 1172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1681685098
transform 1 0 1180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1681685098
transform 1 0 1228 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1681685098
transform 1 0 1244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1681685098
transform 1 0 1236 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_543
timestamp 1681685098
transform 1 0 1236 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1681685098
transform 1 0 1316 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_747
timestamp 1681685098
transform 1 0 1300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1681685098
transform 1 0 1292 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_535
timestamp 1681685098
transform 1 0 1292 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_787
timestamp 1681685098
transform 1 0 1308 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_527
timestamp 1681685098
transform 1 0 1316 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1681685098
transform 1 0 1308 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1681685098
transform 1 0 1332 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_748
timestamp 1681685098
transform 1 0 1332 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_503
timestamp 1681685098
transform 1 0 1348 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1681685098
transform 1 0 1364 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_749
timestamp 1681685098
transform 1 0 1356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1681685098
transform 1 0 1356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1681685098
transform 1 0 1404 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_545
timestamp 1681685098
transform 1 0 1404 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_751
timestamp 1681685098
transform 1 0 1468 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1681685098
transform 1 0 1468 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1681685098
transform 1 0 1500 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1681685098
transform 1 0 1492 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_536
timestamp 1681685098
transform 1 0 1492 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1681685098
transform 1 0 1572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1681685098
transform 1 0 1596 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1681685098
transform 1 0 1588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1681685098
transform 1 0 1684 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_510
timestamp 1681685098
transform 1 0 1700 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1681685098
transform 1 0 1724 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_753
timestamp 1681685098
transform 1 0 1716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1681685098
transform 1 0 1724 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_512
timestamp 1681685098
transform 1 0 1740 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_721
timestamp 1681685098
transform 1 0 1748 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_522
timestamp 1681685098
transform 1 0 1764 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_755
timestamp 1681685098
transform 1 0 1748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1681685098
transform 1 0 1740 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1681685098
transform 1 0 1764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1681685098
transform 1 0 1828 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_523
timestamp 1681685098
transform 1 0 1844 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_756
timestamp 1681685098
transform 1 0 1844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1681685098
transform 1 0 1852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1681685098
transform 1 0 1860 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1681685098
transform 1 0 1876 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1681685098
transform 1 0 1884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1681685098
transform 1 0 1908 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_546
timestamp 1681685098
transform 1 0 1908 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_759
timestamp 1681685098
transform 1 0 1924 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1681685098
transform 1 0 2012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1681685098
transform 1 0 2028 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1681685098
transform 1 0 1932 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1681685098
transform 1 0 1988 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1681685098
transform 1 0 2028 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_537
timestamp 1681685098
transform 1 0 1988 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1681685098
transform 1 0 2036 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1681685098
transform 1 0 2028 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_806
timestamp 1681685098
transform 1 0 2060 0 1 1115
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_18
timestamp 1681685098
transform 1 0 24 0 1 1070
box -10 -3 10 3
use FILL  FILL_676
timestamp 1681685098
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_678
timestamp 1681685098
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_37
timestamp 1681685098
transform 1 0 88 0 -1 1170
box -8 -3 34 105
use FILL  FILL_682
timestamp 1681685098
transform 1 0 120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_684
timestamp 1681685098
transform 1 0 128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_694
timestamp 1681685098
transform 1 0 136 0 -1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_33
timestamp 1681685098
transform -1 0 168 0 -1 1170
box -8 -3 32 105
use XOR2X1  XOR2X1_1
timestamp 1681685098
transform -1 0 224 0 -1 1170
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1681685098
transform 1 0 224 0 -1 1170
box -8 -3 104 105
use FILL  FILL_695
timestamp 1681685098
transform 1 0 320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_696
timestamp 1681685098
transform 1 0 328 0 -1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_2
timestamp 1681685098
transform -1 0 392 0 -1 1170
box -8 -3 64 105
use FILL  FILL_697
timestamp 1681685098
transform 1 0 392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_698
timestamp 1681685098
transform 1 0 400 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1681685098
transform -1 0 504 0 -1 1170
box -8 -3 104 105
use OAI21X1  OAI21X1_39
timestamp 1681685098
transform 1 0 504 0 -1 1170
box -8 -3 34 105
use INVX2  INVX2_36
timestamp 1681685098
transform -1 0 552 0 -1 1170
box -9 -3 26 105
use FILL  FILL_699
timestamp 1681685098
transform 1 0 552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_700
timestamp 1681685098
transform 1 0 560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_701
timestamp 1681685098
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_702
timestamp 1681685098
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_704
timestamp 1681685098
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_706
timestamp 1681685098
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_709
timestamp 1681685098
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1681685098
transform -1 0 640 0 -1 1170
box -8 -3 40 105
use FILL  FILL_710
timestamp 1681685098
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_712
timestamp 1681685098
transform 1 0 648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_714
timestamp 1681685098
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1681685098
transform 1 0 664 0 -1 1170
box -8 -3 104 105
use AOI21X1  AOI21X1_4
timestamp 1681685098
transform 1 0 760 0 -1 1170
box -7 -3 39 105
use INVX2  INVX2_37
timestamp 1681685098
transform -1 0 808 0 -1 1170
box -9 -3 26 105
use FILL  FILL_721
timestamp 1681685098
transform 1 0 808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_722
timestamp 1681685098
transform 1 0 816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_723
timestamp 1681685098
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_725
timestamp 1681685098
transform 1 0 832 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_39
timestamp 1681685098
transform 1 0 840 0 -1 1170
box -9 -3 26 105
use OR2X1  OR2X1_30
timestamp 1681685098
transform -1 0 888 0 -1 1170
box -8 -3 40 105
use FILL  FILL_731
timestamp 1681685098
transform 1 0 888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_733
timestamp 1681685098
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_735
timestamp 1681685098
transform 1 0 904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_737
timestamp 1681685098
transform 1 0 912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_739
timestamp 1681685098
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_741
timestamp 1681685098
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_743
timestamp 1681685098
transform 1 0 936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_744
timestamp 1681685098
transform 1 0 944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_745
timestamp 1681685098
transform 1 0 952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_746
timestamp 1681685098
transform 1 0 960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_747
timestamp 1681685098
transform 1 0 968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_749
timestamp 1681685098
transform 1 0 976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_751
timestamp 1681685098
transform 1 0 984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_753
timestamp 1681685098
transform 1 0 992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_755
timestamp 1681685098
transform 1 0 1000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_759
timestamp 1681685098
transform 1 0 1008 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_40
timestamp 1681685098
transform -1 0 1032 0 -1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_42
timestamp 1681685098
transform -1 0 1064 0 -1 1170
box -8 -3 34 105
use FILL  FILL_760
timestamp 1681685098
transform 1 0 1064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_761
timestamp 1681685098
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_763
timestamp 1681685098
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_765
timestamp 1681685098
transform 1 0 1088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_767
timestamp 1681685098
transform 1 0 1096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_773
timestamp 1681685098
transform 1 0 1104 0 -1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_3
timestamp 1681685098
transform -1 0 1168 0 -1 1170
box -8 -3 64 105
use FILL  FILL_774
timestamp 1681685098
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_4
timestamp 1681685098
transform 1 0 1176 0 -1 1170
box -8 -3 64 105
use FILL  FILL_782
timestamp 1681685098
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use BUFX2  BUFX2_2
timestamp 1681685098
transform -1 0 1264 0 -1 1170
box -5 -3 28 105
use FILL  FILL_783
timestamp 1681685098
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_784
timestamp 1681685098
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_785
timestamp 1681685098
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_786
timestamp 1681685098
transform 1 0 1288 0 -1 1170
box -8 -3 16 105
use AND2X2  AND2X2_4
timestamp 1681685098
transform 1 0 1296 0 -1 1170
box -8 -3 40 105
use FILL  FILL_787
timestamp 1681685098
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_788
timestamp 1681685098
transform 1 0 1336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_789
timestamp 1681685098
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_5
timestamp 1681685098
transform 1 0 1352 0 -1 1170
box -8 -3 64 105
use FILL  FILL_790
timestamp 1681685098
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_792
timestamp 1681685098
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_794
timestamp 1681685098
transform 1 0 1424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_796
timestamp 1681685098
transform 1 0 1432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_804
timestamp 1681685098
transform 1 0 1440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_805
timestamp 1681685098
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_806
timestamp 1681685098
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_807
timestamp 1681685098
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use BUFX2  BUFX2_4
timestamp 1681685098
transform -1 0 1496 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1681685098
transform -1 0 1520 0 -1 1170
box -5 -3 28 105
use FILL  FILL_808
timestamp 1681685098
transform 1 0 1520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_809
timestamp 1681685098
transform 1 0 1528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_810
timestamp 1681685098
transform 1 0 1536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_811
timestamp 1681685098
transform 1 0 1544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_812
timestamp 1681685098
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_813
timestamp 1681685098
transform 1 0 1560 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1681685098
transform -1 0 1592 0 -1 1170
box -8 -3 32 105
use FILL  FILL_814
timestamp 1681685098
transform 1 0 1592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_815
timestamp 1681685098
transform 1 0 1600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_816
timestamp 1681685098
transform 1 0 1608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_818
timestamp 1681685098
transform 1 0 1616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_820
timestamp 1681685098
transform 1 0 1624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_822
timestamp 1681685098
transform 1 0 1632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_825
timestamp 1681685098
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_41
timestamp 1681685098
transform -1 0 1664 0 -1 1170
box -9 -3 26 105
use FILL  FILL_826
timestamp 1681685098
transform 1 0 1664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_827
timestamp 1681685098
transform 1 0 1672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_828
timestamp 1681685098
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_830
timestamp 1681685098
transform 1 0 1688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_832
timestamp 1681685098
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_834
timestamp 1681685098
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_838
timestamp 1681685098
transform 1 0 1712 0 -1 1170
box -8 -3 16 105
use BUFX2  BUFX2_6
timestamp 1681685098
transform -1 0 1744 0 -1 1170
box -5 -3 28 105
use NOR2X1  NOR2X1_13
timestamp 1681685098
transform 1 0 1744 0 -1 1170
box -8 -3 32 105
use FILL  FILL_839
timestamp 1681685098
transform 1 0 1768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_840
timestamp 1681685098
transform 1 0 1776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_841
timestamp 1681685098
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_843
timestamp 1681685098
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_845
timestamp 1681685098
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_850
timestamp 1681685098
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_851
timestamp 1681685098
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_852
timestamp 1681685098
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_42
timestamp 1681685098
transform -1 0 1848 0 -1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_44
timestamp 1681685098
transform 1 0 1848 0 -1 1170
box -8 -3 34 105
use FILL  FILL_853
timestamp 1681685098
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_854
timestamp 1681685098
transform 1 0 1888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_855
timestamp 1681685098
transform 1 0 1896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_856
timestamp 1681685098
transform 1 0 1904 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_43
timestamp 1681685098
transform -1 0 1928 0 -1 1170
box -9 -3 26 105
use M3_M2  M3_M2_548
timestamp 1681685098
transform 1 0 1988 0 1 1075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_41
timestamp 1681685098
transform -1 0 2024 0 -1 1170
box -8 -3 104 105
use NAND2X1  NAND2X1_36
timestamp 1681685098
transform 1 0 2024 0 -1 1170
box -8 -3 32 105
use FILL  FILL_857
timestamp 1681685098
transform 1 0 2048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_859
timestamp 1681685098
transform 1 0 2056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_861
timestamp 1681685098
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_863
timestamp 1681685098
transform 1 0 2072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_865
timestamp 1681685098
transform 1 0 2080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_867
timestamp 1681685098
transform 1 0 2088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_869
timestamp 1681685098
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_871
timestamp 1681685098
transform 1 0 2104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_873
timestamp 1681685098
transform 1 0 2112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_875
timestamp 1681685098
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_877
timestamp 1681685098
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_879
timestamp 1681685098
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_19
timestamp 1681685098
transform 1 0 2194 0 1 1070
box -10 -3 10 3
use M3_M2  M3_M2_559
timestamp 1681685098
transform 1 0 180 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_815
timestamp 1681685098
transform 1 0 180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1681685098
transform 1 0 188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1681685098
transform 1 0 156 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_568
timestamp 1681685098
transform 1 0 228 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_817
timestamp 1681685098
transform 1 0 228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1681685098
transform 1 0 204 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_569
timestamp 1681685098
transform 1 0 252 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_856
timestamp 1681685098
transform 1 0 236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1681685098
transform 1 0 244 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_599
timestamp 1681685098
transform 1 0 244 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1681685098
transform 1 0 284 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1681685098
transform 1 0 308 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1681685098
transform 1 0 324 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_818
timestamp 1681685098
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_573
timestamp 1681685098
transform 1 0 444 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_819
timestamp 1681685098
transform 1 0 324 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1681685098
transform 1 0 340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1681685098
transform 1 0 380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1681685098
transform 1 0 436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1681685098
transform 1 0 308 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1681685098
transform 1 0 316 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_600
timestamp 1681685098
transform 1 0 316 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1681685098
transform 1 0 460 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_860
timestamp 1681685098
transform 1 0 356 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_593
timestamp 1681685098
transform 1 0 436 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_861
timestamp 1681685098
transform 1 0 444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1681685098
transform 1 0 460 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_560
timestamp 1681685098
transform 1 0 484 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_823
timestamp 1681685098
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1681685098
transform 1 0 484 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_601
timestamp 1681685098
transform 1 0 468 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_810
timestamp 1681685098
transform 1 0 492 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_588
timestamp 1681685098
transform 1 0 508 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_864
timestamp 1681685098
transform 1 0 500 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_602
timestamp 1681685098
transform 1 0 500 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1681685098
transform 1 0 492 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1681685098
transform 1 0 540 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_824
timestamp 1681685098
transform 1 0 532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1681685098
transform 1 0 548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1681685098
transform 1 0 540 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_589
timestamp 1681685098
transform 1 0 564 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_883
timestamp 1681685098
transform 1 0 556 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_610
timestamp 1681685098
transform 1 0 548 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_866
timestamp 1681685098
transform 1 0 604 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_575
timestamp 1681685098
transform 1 0 628 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_826
timestamp 1681685098
transform 1 0 628 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_594
timestamp 1681685098
transform 1 0 628 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1681685098
transform 1 0 780 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_827
timestamp 1681685098
transform 1 0 788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1681685098
transform 1 0 748 0 1 1007
box -2 -2 2 2
use M3_M2  M3_M2_603
timestamp 1681685098
transform 1 0 748 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1681685098
transform 1 0 876 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_828
timestamp 1681685098
transform 1 0 868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1681685098
transform 1 0 876 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_549
timestamp 1681685098
transform 1 0 884 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_867
timestamp 1681685098
transform 1 0 884 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_578
timestamp 1681685098
transform 1 0 908 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_868
timestamp 1681685098
transform 1 0 908 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_604
timestamp 1681685098
transform 1 0 908 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1681685098
transform 1 0 924 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_830
timestamp 1681685098
transform 1 0 924 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_590
timestamp 1681685098
transform 1 0 940 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1681685098
transform 1 0 1124 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_831
timestamp 1681685098
transform 1 0 964 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1681685098
transform 1 0 1020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1681685098
transform 1 0 1060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1681685098
transform 1 0 1116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1681685098
transform 1 0 1124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1681685098
transform 1 0 940 0 1 1007
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1681685098
transform 1 0 1036 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_595
timestamp 1681685098
transform 1 0 1116 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1681685098
transform 1 0 1020 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1681685098
transform 1 0 1036 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1681685098
transform 1 0 1148 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1681685098
transform 1 0 1140 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_836
timestamp 1681685098
transform 1 0 1148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1681685098
transform 1 0 1140 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_551
timestamp 1681685098
transform 1 0 1180 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_837
timestamp 1681685098
transform 1 0 1180 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_552
timestamp 1681685098
transform 1 0 1244 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1681685098
transform 1 0 1316 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1681685098
transform 1 0 1284 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1681685098
transform 1 0 1308 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_838
timestamp 1681685098
transform 1 0 1308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1681685098
transform 1 0 1196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1681685098
transform 1 0 1204 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_607
timestamp 1681685098
transform 1 0 1196 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1681685098
transform 1 0 1212 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_884
timestamp 1681685098
transform 1 0 1220 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_562
timestamp 1681685098
transform 1 0 1332 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1681685098
transform 1 0 1356 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1681685098
transform 1 0 1460 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_839
timestamp 1681685098
transform 1 0 1348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1681685098
transform 1 0 1356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1681685098
transform 1 0 1364 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1681685098
transform 1 0 1340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1681685098
transform 1 0 1348 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1681685098
transform 1 0 1460 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1681685098
transform 1 0 1468 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_608
timestamp 1681685098
transform 1 0 1436 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_885
timestamp 1681685098
transform 1 0 1452 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_553
timestamp 1681685098
transform 1 0 1500 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1681685098
transform 1 0 1508 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_842
timestamp 1681685098
transform 1 0 1500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1681685098
transform 1 0 1516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1681685098
transform 1 0 1540 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_611
timestamp 1681685098
transform 1 0 1532 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1681685098
transform 1 0 1588 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1681685098
transform 1 0 1580 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_845
timestamp 1681685098
transform 1 0 1580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1681685098
transform 1 0 1588 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1681685098
transform 1 0 1652 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_550
timestamp 1681685098
transform 1 0 1676 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_811
timestamp 1681685098
transform 1 0 1676 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_565
timestamp 1681685098
transform 1 0 1716 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_846
timestamp 1681685098
transform 1 0 1716 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_554
timestamp 1681685098
transform 1 0 1732 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_807
timestamp 1681685098
transform 1 0 1732 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_566
timestamp 1681685098
transform 1 0 1740 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_808
timestamp 1681685098
transform 1 0 1748 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_585
timestamp 1681685098
transform 1 0 1740 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_847
timestamp 1681685098
transform 1 0 1740 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_567
timestamp 1681685098
transform 1 0 1788 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_812
timestamp 1681685098
transform 1 0 1796 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1681685098
transform 1 0 1788 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_555
timestamp 1681685098
transform 1 0 1844 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_809
timestamp 1681685098
transform 1 0 1836 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1681685098
transform 1 0 1812 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_586
timestamp 1681685098
transform 1 0 1828 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_814
timestamp 1681685098
transform 1 0 1844 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1681685098
transform 1 0 1828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1681685098
transform 1 0 1812 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_592
timestamp 1681685098
transform 1 0 1844 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1681685098
transform 1 0 1988 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_850
timestamp 1681685098
transform 1 0 1972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1681685098
transform 1 0 2028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1681685098
transform 1 0 1948 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_597
timestamp 1681685098
transform 1 0 2028 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_881
timestamp 1681685098
transform 1 0 2036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1681685098
transform 1 0 2036 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_598
timestamp 1681685098
transform 1 0 2052 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1681685098
transform 1 0 2068 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_882
timestamp 1681685098
transform 1 0 2116 0 1 1005
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_20
timestamp 1681685098
transform 1 0 48 0 1 970
box -10 -3 10 3
use FILL  FILL_880
timestamp 1681685098
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_882
timestamp 1681685098
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_884
timestamp 1681685098
transform 1 0 88 0 1 970
box -8 -3 16 105
use FILL  FILL_886
timestamp 1681685098
transform 1 0 96 0 1 970
box -8 -3 16 105
use FILL  FILL_888
timestamp 1681685098
transform 1 0 104 0 1 970
box -8 -3 16 105
use FILL  FILL_890
timestamp 1681685098
transform 1 0 112 0 1 970
box -8 -3 16 105
use FILL  FILL_892
timestamp 1681685098
transform 1 0 120 0 1 970
box -8 -3 16 105
use FILL  FILL_893
timestamp 1681685098
transform 1 0 128 0 1 970
box -8 -3 16 105
use FILL  FILL_894
timestamp 1681685098
transform 1 0 136 0 1 970
box -8 -3 16 105
use FILL  FILL_895
timestamp 1681685098
transform 1 0 144 0 1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_6
timestamp 1681685098
transform 1 0 152 0 1 970
box -8 -3 64 105
use AND2X2  AND2X2_5
timestamp 1681685098
transform -1 0 240 0 1 970
box -8 -3 40 105
use FILL  FILL_896
timestamp 1681685098
transform 1 0 240 0 1 970
box -8 -3 16 105
use FILL  FILL_897
timestamp 1681685098
transform 1 0 248 0 1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_7
timestamp 1681685098
transform 1 0 256 0 1 970
box -8 -3 64 105
use AND2X2  AND2X2_6
timestamp 1681685098
transform 1 0 312 0 1 970
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1681685098
transform 1 0 344 0 1 970
box -8 -3 104 105
use INVX2  INVX2_44
timestamp 1681685098
transform 1 0 440 0 1 970
box -9 -3 26 105
use OAI21X1  OAI21X1_45
timestamp 1681685098
transform 1 0 456 0 1 970
box -8 -3 34 105
use FILL  FILL_898
timestamp 1681685098
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_899
timestamp 1681685098
transform 1 0 496 0 1 970
box -8 -3 16 105
use FILL  FILL_915
timestamp 1681685098
transform 1 0 504 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1681685098
transform -1 0 552 0 1 970
box -8 -3 46 105
use FILL  FILL_916
timestamp 1681685098
transform 1 0 552 0 1 970
box -8 -3 16 105
use FILL  FILL_917
timestamp 1681685098
transform 1 0 560 0 1 970
box -8 -3 16 105
use FILL  FILL_918
timestamp 1681685098
transform 1 0 568 0 1 970
box -8 -3 16 105
use FILL  FILL_919
timestamp 1681685098
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_920
timestamp 1681685098
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_925
timestamp 1681685098
transform 1 0 592 0 1 970
box -8 -3 16 105
use FILL  FILL_927
timestamp 1681685098
transform 1 0 600 0 1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_14
timestamp 1681685098
transform 1 0 608 0 1 970
box -8 -3 32 105
use FILL  FILL_929
timestamp 1681685098
transform 1 0 632 0 1 970
box -8 -3 16 105
use FILL  FILL_930
timestamp 1681685098
transform 1 0 640 0 1 970
box -8 -3 16 105
use FILL  FILL_932
timestamp 1681685098
transform 1 0 648 0 1 970
box -8 -3 16 105
use FILL  FILL_934
timestamp 1681685098
transform 1 0 656 0 1 970
box -8 -3 16 105
use FILL  FILL_936
timestamp 1681685098
transform 1 0 664 0 1 970
box -8 -3 16 105
use FILL  FILL_937
timestamp 1681685098
transform 1 0 672 0 1 970
box -8 -3 16 105
use FILL  FILL_938
timestamp 1681685098
transform 1 0 680 0 1 970
box -8 -3 16 105
use FILL  FILL_939
timestamp 1681685098
transform 1 0 688 0 1 970
box -8 -3 16 105
use FILL  FILL_940
timestamp 1681685098
transform 1 0 696 0 1 970
box -8 -3 16 105
use FILL  FILL_941
timestamp 1681685098
transform 1 0 704 0 1 970
box -8 -3 16 105
use FILL  FILL_944
timestamp 1681685098
transform 1 0 712 0 1 970
box -8 -3 16 105
use FILL  FILL_946
timestamp 1681685098
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_948
timestamp 1681685098
transform 1 0 728 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1681685098
transform 1 0 736 0 1 970
box -8 -3 104 105
use FILL  FILL_950
timestamp 1681685098
transform 1 0 832 0 1 970
box -8 -3 16 105
use FILL  FILL_956
timestamp 1681685098
transform 1 0 840 0 1 970
box -8 -3 16 105
use FILL  FILL_958
timestamp 1681685098
transform 1 0 848 0 1 970
box -8 -3 16 105
use FILL  FILL_960
timestamp 1681685098
transform 1 0 856 0 1 970
box -8 -3 16 105
use FILL  FILL_962
timestamp 1681685098
transform 1 0 864 0 1 970
box -8 -3 16 105
use FILL  FILL_963
timestamp 1681685098
transform 1 0 872 0 1 970
box -8 -3 16 105
use FILL  FILL_964
timestamp 1681685098
transform 1 0 880 0 1 970
box -8 -3 16 105
use INVX2  INVX2_47
timestamp 1681685098
transform 1 0 888 0 1 970
box -9 -3 26 105
use BUFX2  BUFX2_7
timestamp 1681685098
transform -1 0 928 0 1 970
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1681685098
transform 1 0 928 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1681685098
transform 1 0 1024 0 1 970
box -8 -3 104 105
use BUFX2  BUFX2_8
timestamp 1681685098
transform 1 0 1120 0 1 970
box -5 -3 28 105
use FILL  FILL_966
timestamp 1681685098
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_992
timestamp 1681685098
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_994
timestamp 1681685098
transform 1 0 1160 0 1 970
box -8 -3 16 105
use FILL  FILL_995
timestamp 1681685098
transform 1 0 1168 0 1 970
box -8 -3 16 105
use BUFX2  BUFX2_9
timestamp 1681685098
transform 1 0 1176 0 1 970
box -5 -3 28 105
use FILL  FILL_996
timestamp 1681685098
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FAX1  FAX1_1
timestamp 1681685098
transform -1 0 1328 0 1 970
box -5 -3 126 105
use FILL  FILL_997
timestamp 1681685098
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_998
timestamp 1681685098
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FAX1  FAX1_2
timestamp 1681685098
transform 1 0 1344 0 1 970
box -5 -3 126 105
use FILL  FILL_999
timestamp 1681685098
transform 1 0 1464 0 1 970
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1681685098
transform 1 0 1472 0 1 970
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1681685098
transform 1 0 1480 0 1 970
box -8 -3 16 105
use AND2X2  AND2X2_13
timestamp 1681685098
transform 1 0 1488 0 1 970
box -8 -3 40 105
use FILL  FILL_1013
timestamp 1681685098
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1681685098
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1681685098
transform 1 0 1536 0 1 970
box -8 -3 16 105
use INVX2  INVX2_49
timestamp 1681685098
transform -1 0 1560 0 1 970
box -9 -3 26 105
use AND2X2  AND2X2_14
timestamp 1681685098
transform -1 0 1592 0 1 970
box -8 -3 40 105
use FILL  FILL_1021
timestamp 1681685098
transform 1 0 1592 0 1 970
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1681685098
transform 1 0 1600 0 1 970
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1681685098
transform 1 0 1608 0 1 970
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1681685098
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1681685098
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1681685098
transform 1 0 1632 0 1 970
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1681685098
transform 1 0 1640 0 1 970
box -8 -3 16 105
use BUFX2  BUFX2_10
timestamp 1681685098
transform -1 0 1672 0 1 970
box -5 -3 28 105
use FILL  FILL_1028
timestamp 1681685098
transform 1 0 1672 0 1 970
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1681685098
transform 1 0 1680 0 1 970
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1681685098
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1681685098
transform 1 0 1696 0 1 970
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1681685098
transform 1 0 1704 0 1 970
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1681685098
transform 1 0 1712 0 1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_12
timestamp 1681685098
transform -1 0 1752 0 1 970
box -8 -3 40 105
use FILL  FILL_1037
timestamp 1681685098
transform 1 0 1752 0 1 970
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1681685098
transform 1 0 1760 0 1 970
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1681685098
transform 1 0 1768 0 1 970
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1681685098
transform 1 0 1776 0 1 970
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1681685098
transform 1 0 1784 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_37
timestamp 1681685098
transform -1 0 1816 0 1 970
box -8 -3 32 105
use NAND3X1  NAND3X1_13
timestamp 1681685098
transform 1 0 1816 0 1 970
box -8 -3 40 105
use FILL  FILL_1051
timestamp 1681685098
transform 1 0 1848 0 1 970
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1681685098
transform 1 0 1856 0 1 970
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1681685098
transform 1 0 1864 0 1 970
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1681685098
transform 1 0 1872 0 1 970
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1681685098
transform 1 0 1880 0 1 970
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1681685098
transform 1 0 1888 0 1 970
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1681685098
transform 1 0 1896 0 1 970
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1681685098
transform 1 0 1904 0 1 970
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1681685098
transform 1 0 1912 0 1 970
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1681685098
transform 1 0 1920 0 1 970
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1681685098
transform 1 0 1928 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1681685098
transform 1 0 1936 0 1 970
box -8 -3 104 105
use NOR2X1  NOR2X1_15
timestamp 1681685098
transform 1 0 2032 0 1 970
box -8 -3 32 105
use FILL  FILL_1062
timestamp 1681685098
transform 1 0 2056 0 1 970
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1681685098
transform 1 0 2064 0 1 970
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1681685098
transform 1 0 2072 0 1 970
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1681685098
transform 1 0 2080 0 1 970
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1681685098
transform 1 0 2088 0 1 970
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1681685098
transform 1 0 2096 0 1 970
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1681685098
transform 1 0 2104 0 1 970
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1681685098
transform 1 0 2112 0 1 970
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1681685098
transform 1 0 2120 0 1 970
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1681685098
transform 1 0 2128 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_613
timestamp 1681685098
transform 1 0 2148 0 1 975
box -3 -3 3 3
use FILL  FILL_1072
timestamp 1681685098
transform 1 0 2136 0 1 970
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_21
timestamp 1681685098
transform 1 0 2170 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_624
timestamp 1681685098
transform 1 0 124 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_890
timestamp 1681685098
transform 1 0 124 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_625
timestamp 1681685098
transform 1 0 180 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_891
timestamp 1681685098
transform 1 0 172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1681685098
transform 1 0 180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1681685098
transform 1 0 156 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_618
timestamp 1681685098
transform 1 0 212 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1681685098
transform 1 0 236 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_893
timestamp 1681685098
transform 1 0 212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1681685098
transform 1 0 260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1681685098
transform 1 0 268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1681685098
transform 1 0 188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1681685098
transform 1 0 204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1681685098
transform 1 0 236 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_647
timestamp 1681685098
transform 1 0 172 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1681685098
transform 1 0 188 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1681685098
transform 1 0 156 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1681685098
transform 1 0 236 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_896
timestamp 1681685098
transform 1 0 324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1681685098
transform 1 0 300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1681685098
transform 1 0 316 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_650
timestamp 1681685098
transform 1 0 300 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1681685098
transform 1 0 324 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1681685098
transform 1 0 364 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_897
timestamp 1681685098
transform 1 0 364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1681685098
transform 1 0 380 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1681685098
transform 1 0 380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1681685098
transform 1 0 396 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1681685098
transform 1 0 380 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_620
timestamp 1681685098
transform 1 0 444 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1681685098
transform 1 0 436 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_899
timestamp 1681685098
transform 1 0 428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1681685098
transform 1 0 420 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_659
timestamp 1681685098
transform 1 0 420 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1681685098
transform 1 0 460 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_900
timestamp 1681685098
transform 1 0 460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1681685098
transform 1 0 468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1681685098
transform 1 0 484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1681685098
transform 1 0 476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1681685098
transform 1 0 492 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_660
timestamp 1681685098
transform 1 0 492 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1681685098
transform 1 0 476 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1681685098
transform 1 0 556 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_903
timestamp 1681685098
transform 1 0 532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1681685098
transform 1 0 524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1681685098
transform 1 0 580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1681685098
transform 1 0 604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1681685098
transform 1 0 620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1681685098
transform 1 0 668 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1681685098
transform 1 0 676 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_642
timestamp 1681685098
transform 1 0 684 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_952
timestamp 1681685098
transform 1 0 692 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_668
timestamp 1681685098
transform 1 0 692 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_906
timestamp 1681685098
transform 1 0 732 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_633
timestamp 1681685098
transform 1 0 740 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1681685098
transform 1 0 732 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1681685098
transform 1 0 772 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_907
timestamp 1681685098
transform 1 0 780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1681685098
transform 1 0 788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1681685098
transform 1 0 756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1681685098
transform 1 0 772 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_643
timestamp 1681685098
transform 1 0 780 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1681685098
transform 1 0 756 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_983
timestamp 1681685098
transform 1 0 788 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_629
timestamp 1681685098
transform 1 0 812 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_909
timestamp 1681685098
transform 1 0 812 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_644
timestamp 1681685098
transform 1 0 812 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1681685098
transform 1 0 796 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_910
timestamp 1681685098
transform 1 0 836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1681685098
transform 1 0 868 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_653
timestamp 1681685098
transform 1 0 868 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_912
timestamp 1681685098
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1681685098
transform 1 0 980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1681685098
transform 1 0 972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1681685098
transform 1 0 980 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_630
timestamp 1681685098
transform 1 0 1028 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_914
timestamp 1681685098
transform 1 0 1028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1681685098
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1681685098
transform 1 0 1060 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1681685098
transform 1 0 1060 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_654
timestamp 1681685098
transform 1 0 1060 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_984
timestamp 1681685098
transform 1 0 1068 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_661
timestamp 1681685098
transform 1 0 1068 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_916
timestamp 1681685098
transform 1 0 1172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1681685098
transform 1 0 1188 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_645
timestamp 1681685098
transform 1 0 1172 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_959
timestamp 1681685098
transform 1 0 1180 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_662
timestamp 1681685098
transform 1 0 1180 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_918
timestamp 1681685098
transform 1 0 1212 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_669
timestamp 1681685098
transform 1 0 1212 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1681685098
transform 1 0 1260 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_919
timestamp 1681685098
transform 1 0 1252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1681685098
transform 1 0 1260 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_632
timestamp 1681685098
transform 1 0 1316 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_921
timestamp 1681685098
transform 1 0 1316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1681685098
transform 1 0 1260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1681685098
transform 1 0 1284 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_646
timestamp 1681685098
transform 1 0 1292 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_962
timestamp 1681685098
transform 1 0 1308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1681685098
transform 1 0 1324 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_655
timestamp 1681685098
transform 1 0 1260 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1681685098
transform 1 0 1284 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1681685098
transform 1 0 1324 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1681685098
transform 1 0 1348 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_922
timestamp 1681685098
transform 1 0 1436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1681685098
transform 1 0 1348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1681685098
transform 1 0 1356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1681685098
transform 1 0 1412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1681685098
transform 1 0 1452 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_665
timestamp 1681685098
transform 1 0 1356 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_968
timestamp 1681685098
transform 1 0 1492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1681685098
transform 1 0 1516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1681685098
transform 1 0 1516 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_666
timestamp 1681685098
transform 1 0 1516 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_887
timestamp 1681685098
transform 1 0 1636 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1681685098
transform 1 0 1532 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_636
timestamp 1681685098
transform 1 0 1548 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1681685098
transform 1 0 1636 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_925
timestamp 1681685098
transform 1 0 1644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1681685098
transform 1 0 1548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1681685098
transform 1 0 1668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1681685098
transform 1 0 1684 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_638
timestamp 1681685098
transform 1 0 1692 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_971
timestamp 1681685098
transform 1 0 1660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1681685098
transform 1 0 1676 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1681685098
transform 1 0 1692 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_670
timestamp 1681685098
transform 1 0 1652 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1681685098
transform 1 0 1684 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_928
timestamp 1681685098
transform 1 0 1756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1681685098
transform 1 0 1788 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1681685098
transform 1 0 1820 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1681685098
transform 1 0 1836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1681685098
transform 1 0 1812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1681685098
transform 1 0 1820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1681685098
transform 1 0 1804 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_639
timestamp 1681685098
transform 1 0 1908 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_931
timestamp 1681685098
transform 1 0 1932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1681685098
transform 1 0 1908 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_672
timestamp 1681685098
transform 1 0 1900 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1681685098
transform 1 0 1932 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1681685098
transform 1 0 1956 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_888
timestamp 1681685098
transform 1 0 1956 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1681685098
transform 1 0 1956 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_615
timestamp 1681685098
transform 1 0 1988 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1681685098
transform 1 0 1980 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_889
timestamp 1681685098
transform 1 0 1988 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_616
timestamp 1681685098
transform 1 0 2012 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1681685098
transform 1 0 2036 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_932
timestamp 1681685098
transform 1 0 1980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1681685098
transform 1 0 1996 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1681685098
transform 1 0 1980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1681685098
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_640
timestamp 1681685098
transform 1 0 2052 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1681685098
transform 1 0 2068 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1681685098
transform 1 0 2140 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_935
timestamp 1681685098
transform 1 0 2116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1681685098
transform 1 0 2140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1681685098
transform 1 0 2012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1681685098
transform 1 0 2052 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1681685098
transform 1 0 2148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1681685098
transform 1 0 2116 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_674
timestamp 1681685098
transform 1 0 2028 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1681685098
transform 1 0 2116 0 1 885
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_22
timestamp 1681685098
transform 1 0 24 0 1 870
box -10 -3 10 3
use FILL  FILL_881
timestamp 1681685098
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_883
timestamp 1681685098
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_885
timestamp 1681685098
transform 1 0 88 0 -1 970
box -8 -3 16 105
use FILL  FILL_887
timestamp 1681685098
transform 1 0 96 0 -1 970
box -8 -3 16 105
use FILL  FILL_889
timestamp 1681685098
transform 1 0 104 0 -1 970
box -8 -3 16 105
use FILL  FILL_891
timestamp 1681685098
transform 1 0 112 0 -1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_8
timestamp 1681685098
transform 1 0 120 0 -1 970
box -8 -3 64 105
use AND2X2  AND2X2_7
timestamp 1681685098
transform 1 0 176 0 -1 970
box -8 -3 40 105
use XOR2X1  XOR2X1_9
timestamp 1681685098
transform 1 0 208 0 -1 970
box -8 -3 64 105
use FILL  FILL_900
timestamp 1681685098
transform 1 0 264 0 -1 970
box -8 -3 16 105
use FILL  FILL_901
timestamp 1681685098
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_902
timestamp 1681685098
transform 1 0 280 0 -1 970
box -8 -3 16 105
use AND2X2  AND2X2_8
timestamp 1681685098
transform 1 0 288 0 -1 970
box -8 -3 40 105
use FILL  FILL_903
timestamp 1681685098
transform 1 0 320 0 -1 970
box -8 -3 16 105
use FILL  FILL_904
timestamp 1681685098
transform 1 0 328 0 -1 970
box -8 -3 16 105
use FILL  FILL_905
timestamp 1681685098
transform 1 0 336 0 -1 970
box -8 -3 16 105
use FILL  FILL_906
timestamp 1681685098
transform 1 0 344 0 -1 970
box -8 -3 16 105
use FILL  FILL_907
timestamp 1681685098
transform 1 0 352 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_45
timestamp 1681685098
transform 1 0 360 0 -1 970
box -9 -3 26 105
use OAI21X1  OAI21X1_46
timestamp 1681685098
transform -1 0 408 0 -1 970
box -8 -3 34 105
use FILL  FILL_908
timestamp 1681685098
transform 1 0 408 0 -1 970
box -8 -3 16 105
use FILL  FILL_909
timestamp 1681685098
transform 1 0 416 0 -1 970
box -8 -3 16 105
use FILL  FILL_910
timestamp 1681685098
transform 1 0 424 0 -1 970
box -8 -3 16 105
use FILL  FILL_911
timestamp 1681685098
transform 1 0 432 0 -1 970
box -8 -3 16 105
use FILL  FILL_912
timestamp 1681685098
transform 1 0 440 0 -1 970
box -8 -3 16 105
use FILL  FILL_913
timestamp 1681685098
transform 1 0 448 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_0
timestamp 1681685098
transform -1 0 496 0 -1 970
box -8 -3 46 105
use FILL  FILL_914
timestamp 1681685098
transform 1 0 496 0 -1 970
box -8 -3 16 105
use FILL  FILL_921
timestamp 1681685098
transform 1 0 504 0 -1 970
box -8 -3 16 105
use FILL  FILL_922
timestamp 1681685098
transform 1 0 512 0 -1 970
box -8 -3 16 105
use FILL  FILL_923
timestamp 1681685098
transform 1 0 520 0 -1 970
box -8 -3 16 105
use XNOR2X1  XNOR2X1_32
timestamp 1681685098
transform -1 0 584 0 -1 970
box -8 -3 64 105
use FILL  FILL_924
timestamp 1681685098
transform 1 0 584 0 -1 970
box -8 -3 16 105
use FILL  FILL_926
timestamp 1681685098
transform 1 0 592 0 -1 970
box -8 -3 16 105
use FILL  FILL_928
timestamp 1681685098
transform 1 0 600 0 -1 970
box -8 -3 16 105
use AND2X2  AND2X2_9
timestamp 1681685098
transform 1 0 608 0 -1 970
box -8 -3 40 105
use FILL  FILL_931
timestamp 1681685098
transform 1 0 640 0 -1 970
box -8 -3 16 105
use FILL  FILL_933
timestamp 1681685098
transform 1 0 648 0 -1 970
box -8 -3 16 105
use FILL  FILL_935
timestamp 1681685098
transform 1 0 656 0 -1 970
box -8 -3 16 105
use FILL  FILL_942
timestamp 1681685098
transform 1 0 664 0 -1 970
box -8 -3 16 105
use AND2X2  AND2X2_10
timestamp 1681685098
transform -1 0 704 0 -1 970
box -8 -3 40 105
use FILL  FILL_943
timestamp 1681685098
transform 1 0 704 0 -1 970
box -8 -3 16 105
use FILL  FILL_945
timestamp 1681685098
transform 1 0 712 0 -1 970
box -8 -3 16 105
use FILL  FILL_947
timestamp 1681685098
transform 1 0 720 0 -1 970
box -8 -3 16 105
use FILL  FILL_949
timestamp 1681685098
transform 1 0 728 0 -1 970
box -8 -3 16 105
use FILL  FILL_951
timestamp 1681685098
transform 1 0 736 0 -1 970
box -8 -3 16 105
use FILL  FILL_952
timestamp 1681685098
transform 1 0 744 0 -1 970
box -8 -3 16 105
use AND2X2  AND2X2_11
timestamp 1681685098
transform -1 0 784 0 -1 970
box -8 -3 40 105
use OAI21X1  OAI21X1_47
timestamp 1681685098
transform -1 0 816 0 -1 970
box -8 -3 34 105
use FILL  FILL_953
timestamp 1681685098
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_954
timestamp 1681685098
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_955
timestamp 1681685098
transform 1 0 832 0 -1 970
box -8 -3 16 105
use FILL  FILL_957
timestamp 1681685098
transform 1 0 840 0 -1 970
box -8 -3 16 105
use FILL  FILL_959
timestamp 1681685098
transform 1 0 848 0 -1 970
box -8 -3 16 105
use FILL  FILL_961
timestamp 1681685098
transform 1 0 856 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_46
timestamp 1681685098
transform 1 0 864 0 -1 970
box -9 -3 26 105
use FILL  FILL_965
timestamp 1681685098
transform 1 0 880 0 -1 970
box -8 -3 16 105
use FILL  FILL_967
timestamp 1681685098
transform 1 0 888 0 -1 970
box -8 -3 16 105
use FILL  FILL_968
timestamp 1681685098
transform 1 0 896 0 -1 970
box -8 -3 16 105
use FILL  FILL_969
timestamp 1681685098
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_970
timestamp 1681685098
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_971
timestamp 1681685098
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_972
timestamp 1681685098
transform 1 0 928 0 -1 970
box -8 -3 16 105
use FILL  FILL_973
timestamp 1681685098
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_974
timestamp 1681685098
transform 1 0 944 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_48
timestamp 1681685098
transform -1 0 984 0 -1 970
box -8 -3 34 105
use FILL  FILL_975
timestamp 1681685098
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_976
timestamp 1681685098
transform 1 0 992 0 -1 970
box -8 -3 16 105
use FILL  FILL_977
timestamp 1681685098
transform 1 0 1000 0 -1 970
box -8 -3 16 105
use FILL  FILL_978
timestamp 1681685098
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use FILL  FILL_979
timestamp 1681685098
transform 1 0 1016 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_49
timestamp 1681685098
transform 1 0 1024 0 -1 970
box -8 -3 34 105
use FILL  FILL_980
timestamp 1681685098
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use FILL  FILL_981
timestamp 1681685098
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_982
timestamp 1681685098
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_983
timestamp 1681685098
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use FILL  FILL_984
timestamp 1681685098
transform 1 0 1088 0 -1 970
box -8 -3 16 105
use FILL  FILL_985
timestamp 1681685098
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use FILL  FILL_986
timestamp 1681685098
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use FILL  FILL_987
timestamp 1681685098
transform 1 0 1112 0 -1 970
box -8 -3 16 105
use FILL  FILL_988
timestamp 1681685098
transform 1 0 1120 0 -1 970
box -8 -3 16 105
use FILL  FILL_989
timestamp 1681685098
transform 1 0 1128 0 -1 970
box -8 -3 16 105
use FILL  FILL_990
timestamp 1681685098
transform 1 0 1136 0 -1 970
box -8 -3 16 105
use FILL  FILL_991
timestamp 1681685098
transform 1 0 1144 0 -1 970
box -8 -3 16 105
use FILL  FILL_993
timestamp 1681685098
transform 1 0 1152 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_2
timestamp 1681685098
transform 1 0 1160 0 -1 970
box -8 -3 46 105
use FILL  FILL_1000
timestamp 1681685098
transform 1 0 1200 0 -1 970
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1681685098
transform 1 0 1208 0 -1 970
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1681685098
transform 1 0 1216 0 -1 970
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1681685098
transform 1 0 1224 0 -1 970
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1681685098
transform 1 0 1232 0 -1 970
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1681685098
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1681685098
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use XOR2X1  XOR2X1_10
timestamp 1681685098
transform 1 0 1256 0 -1 970
box -8 -3 64 105
use AND2X2  AND2X2_12
timestamp 1681685098
transform 1 0 1312 0 -1 970
box -8 -3 40 105
use FILL  FILL_1007
timestamp 1681685098
transform 1 0 1344 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_676
timestamp 1681685098
transform 1 0 1412 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_46
timestamp 1681685098
transform -1 0 1448 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_48
timestamp 1681685098
transform -1 0 1464 0 -1 970
box -9 -3 26 105
use FILL  FILL_1008
timestamp 1681685098
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1681685098
transform 1 0 1472 0 -1 970
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1681685098
transform 1 0 1480 0 -1 970
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1681685098
transform 1 0 1488 0 -1 970
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1681685098
transform 1 0 1496 0 -1 970
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1681685098
transform 1 0 1504 0 -1 970
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1681685098
transform 1 0 1512 0 -1 970
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1681685098
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_677
timestamp 1681685098
transform 1 0 1588 0 1 875
box -3 -3 3 3
use FAX1  FAX1_3
timestamp 1681685098
transform 1 0 1528 0 -1 970
box -5 -3 126 105
use FILL  FILL_1032
timestamp 1681685098
transform 1 0 1648 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_3
timestamp 1681685098
transform 1 0 1656 0 -1 970
box -8 -3 46 105
use FILL  FILL_1033
timestamp 1681685098
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1681685098
transform 1 0 1704 0 -1 970
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1681685098
transform 1 0 1712 0 -1 970
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1681685098
transform 1 0 1720 0 -1 970
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1681685098
transform 1 0 1728 0 -1 970
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1681685098
transform 1 0 1736 0 -1 970
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1681685098
transform 1 0 1744 0 -1 970
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1681685098
transform 1 0 1752 0 -1 970
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1681685098
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1681685098
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1681685098
transform 1 0 1776 0 -1 970
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1681685098
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1681685098
transform 1 0 1792 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_38
timestamp 1681685098
transform -1 0 1824 0 -1 970
box -8 -3 32 105
use INVX2  INVX2_50
timestamp 1681685098
transform -1 0 1840 0 -1 970
box -9 -3 26 105
use FILL  FILL_1075
timestamp 1681685098
transform 1 0 1840 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1681685098
transform -1 0 1944 0 -1 970
box -8 -3 104 105
use FILL  FILL_1076
timestamp 1681685098
transform 1 0 1944 0 -1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_5
timestamp 1681685098
transform -1 0 1984 0 -1 970
box -7 -3 39 105
use OR2X1  OR2X1_34
timestamp 1681685098
transform 1 0 1984 0 -1 970
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1681685098
transform 1 0 2016 0 -1 970
box -8 -3 104 105
use OAI21X1  OAI21X1_50
timestamp 1681685098
transform -1 0 2144 0 -1 970
box -8 -3 34 105
use top_module_VIA0  top_module_VIA0_23
timestamp 1681685098
transform 1 0 2194 0 1 870
box -10 -3 10 3
use M2_M1  M2_M1_1041
timestamp 1681685098
transform 1 0 84 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1681685098
transform 1 0 100 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_688
timestamp 1681685098
transform 1 0 212 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1681685098
transform 1 0 188 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1681685098
transform 1 0 236 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1681685098
transform 1 0 228 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1681685098
transform 1 0 204 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1681685098
transform 1 0 220 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_995
timestamp 1681685098
transform 1 0 188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1681685098
transform 1 0 156 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_731
timestamp 1681685098
transform 1 0 156 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_996
timestamp 1681685098
transform 1 0 220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1681685098
transform 1 0 236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1681685098
transform 1 0 204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1681685098
transform 1 0 212 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_732
timestamp 1681685098
transform 1 0 212 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1681685098
transform 1 0 260 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1681685098
transform 1 0 292 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_998
timestamp 1681685098
transform 1 0 292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1681685098
transform 1 0 300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1681685098
transform 1 0 268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1681685098
transform 1 0 324 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_722
timestamp 1681685098
transform 1 0 324 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1681685098
transform 1 0 356 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_1046
timestamp 1681685098
transform 1 0 372 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_681
timestamp 1681685098
transform 1 0 388 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1681685098
transform 1 0 412 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1001
timestamp 1681685098
transform 1 0 396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1681685098
transform 1 0 412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1681685098
transform 1 0 388 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_734
timestamp 1681685098
transform 1 0 388 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1681685098
transform 1 0 452 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_1048
timestamp 1681685098
transform 1 0 436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1681685098
transform 1 0 444 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_683
timestamp 1681685098
transform 1 0 468 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1681685098
transform 1 0 492 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1003
timestamp 1681685098
transform 1 0 476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1681685098
transform 1 0 460 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_742
timestamp 1681685098
transform 1 0 460 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_1051
timestamp 1681685098
transform 1 0 508 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1681685098
transform 1 0 516 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_743
timestamp 1681685098
transform 1 0 516 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_1004
timestamp 1681685098
transform 1 0 540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1681685098
transform 1 0 548 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1681685098
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1681685098
transform 1 0 604 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_723
timestamp 1681685098
transform 1 0 604 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1052
timestamp 1681685098
transform 1 0 612 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1681685098
transform 1 0 644 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_724
timestamp 1681685098
transform 1 0 636 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1081
timestamp 1681685098
transform 1 0 628 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1681685098
transform 1 0 652 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1681685098
transform 1 0 668 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1681685098
transform 1 0 668 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_717
timestamp 1681685098
transform 1 0 684 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1008
timestamp 1681685098
transform 1 0 692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1681685098
transform 1 0 740 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1681685098
transform 1 0 772 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_690
timestamp 1681685098
transform 1 0 796 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1681685098
transform 1 0 788 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1010
timestamp 1681685098
transform 1 0 788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1681685098
transform 1 0 796 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_684
timestamp 1681685098
transform 1 0 828 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1681685098
transform 1 0 852 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_1011
timestamp 1681685098
transform 1 0 836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1681685098
transform 1 0 852 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1681685098
transform 1 0 868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1681685098
transform 1 0 828 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_725
timestamp 1681685098
transform 1 0 836 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1681685098
transform 1 0 852 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1056
timestamp 1681685098
transform 1 0 860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1681685098
transform 1 0 956 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_707
timestamp 1681685098
transform 1 0 972 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1014
timestamp 1681685098
transform 1 0 964 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1681685098
transform 1 0 972 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_727
timestamp 1681685098
transform 1 0 964 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1016
timestamp 1681685098
transform 1 0 1004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1681685098
transform 1 0 980 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_728
timestamp 1681685098
transform 1 0 996 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1082
timestamp 1681685098
transform 1 0 996 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1681685098
transform 1 0 1036 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_708
timestamp 1681685098
transform 1 0 1092 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1018
timestamp 1681685098
transform 1 0 1092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1681685098
transform 1 0 1116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1681685098
transform 1 0 1092 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_735
timestamp 1681685098
transform 1 0 1092 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1681685098
transform 1 0 1140 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_1060
timestamp 1681685098
transform 1 0 1132 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_709
timestamp 1681685098
transform 1 0 1156 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1061
timestamp 1681685098
transform 1 0 1156 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_685
timestamp 1681685098
transform 1 0 1188 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1681685098
transform 1 0 1196 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1020
timestamp 1681685098
transform 1 0 1196 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_691
timestamp 1681685098
transform 1 0 1212 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_1021
timestamp 1681685098
transform 1 0 1212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1681685098
transform 1 0 1228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1681685098
transform 1 0 1204 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_692
timestamp 1681685098
transform 1 0 1292 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1681685098
transform 1 0 1260 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1681685098
transform 1 0 1316 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1023
timestamp 1681685098
transform 1 0 1260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1681685098
transform 1 0 1292 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_736
timestamp 1681685098
transform 1 0 1252 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_1063
timestamp 1681685098
transform 1 0 1308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1681685098
transform 1 0 1316 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_737
timestamp 1681685098
transform 1 0 1308 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_1083
timestamp 1681685098
transform 1 0 1316 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_713
timestamp 1681685098
transform 1 0 1340 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1025
timestamp 1681685098
transform 1 0 1340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1681685098
transform 1 0 1356 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_686
timestamp 1681685098
transform 1 0 1380 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1681685098
transform 1 0 1452 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1681685098
transform 1 0 1460 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1681685098
transform 1 0 1388 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_1027
timestamp 1681685098
transform 1 0 1380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1681685098
transform 1 0 1388 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_718
timestamp 1681685098
transform 1 0 1420 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1681685098
transform 1 0 1412 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1681685098
transform 1 0 1476 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_1065
timestamp 1681685098
transform 1 0 1484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1681685098
transform 1 0 1476 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_744
timestamp 1681685098
transform 1 0 1476 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_1029
timestamp 1681685098
transform 1 0 1516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1681685098
transform 1 0 1524 0 1 807
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1681685098
transform 1 0 1540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1681685098
transform 1 0 1556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1681685098
transform 1 0 1588 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_693
timestamp 1681685098
transform 1 0 1620 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1681685098
transform 1 0 1644 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_991
timestamp 1681685098
transform 1 0 1644 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1681685098
transform 1 0 1644 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_703
timestamp 1681685098
transform 1 0 1676 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1681685098
transform 1 0 1668 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_1031
timestamp 1681685098
transform 1 0 1716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1681685098
transform 1 0 1740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1681685098
transform 1 0 1732 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1681685098
transform 1 0 1748 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_679
timestamp 1681685098
transform 1 0 1780 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_1071
timestamp 1681685098
transform 1 0 1788 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1681685098
transform 1 0 1804 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_738
timestamp 1681685098
transform 1 0 1804 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_992
timestamp 1681685098
transform 1 0 1820 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1681685098
transform 1 0 1820 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_719
timestamp 1681685098
transform 1 0 1852 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1073
timestamp 1681685098
transform 1 0 1844 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_739
timestamp 1681685098
transform 1 0 1844 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_1034
timestamp 1681685098
transform 1 0 1924 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1681685098
transform 1 0 1948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1681685098
transform 1 0 1900 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_740
timestamp 1681685098
transform 1 0 1900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1681685098
transform 1 0 1996 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_1036
timestamp 1681685098
transform 1 0 1996 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1681685098
transform 1 0 1988 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_680
timestamp 1681685098
transform 1 0 2028 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1681685098
transform 1 0 2020 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1681685098
transform 1 0 2012 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_1037
timestamp 1681685098
transform 1 0 2020 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1681685098
transform 1 0 2028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1681685098
transform 1 0 2012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1681685098
transform 1 0 1996 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_741
timestamp 1681685098
transform 1 0 2004 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1681685098
transform 1 0 2060 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_993
timestamp 1681685098
transform 1 0 2068 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1681685098
transform 1 0 2060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1681685098
transform 1 0 2052 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1681685098
transform 1 0 2124 0 1 805
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_24
timestamp 1681685098
transform 1 0 48 0 1 770
box -10 -3 10 3
use FILL  FILL_1077
timestamp 1681685098
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1681685098
transform 1 0 80 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_15
timestamp 1681685098
transform 1 0 88 0 1 770
box -8 -3 40 105
use FILL  FILL_1080
timestamp 1681685098
transform 1 0 120 0 1 770
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1681685098
transform 1 0 128 0 1 770
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1681685098
transform 1 0 136 0 1 770
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1681685098
transform 1 0 144 0 1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_12
timestamp 1681685098
transform 1 0 152 0 1 770
box -8 -3 64 105
use AND2X2  AND2X2_16
timestamp 1681685098
transform 1 0 208 0 1 770
box -8 -3 40 105
use FILL  FILL_1085
timestamp 1681685098
transform 1 0 240 0 1 770
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1681685098
transform 1 0 248 0 1 770
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1681685098
transform 1 0 256 0 1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_14
timestamp 1681685098
transform 1 0 264 0 1 770
box -8 -3 64 105
use FILL  FILL_1092
timestamp 1681685098
transform 1 0 320 0 1 770
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1681685098
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1681685098
transform 1 0 336 0 1 770
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1681685098
transform 1 0 344 0 1 770
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1681685098
transform 1 0 352 0 1 770
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1681685098
transform 1 0 360 0 1 770
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1681685098
transform 1 0 368 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_4
timestamp 1681685098
transform -1 0 416 0 1 770
box -8 -3 46 105
use FILL  FILL_1099
timestamp 1681685098
transform 1 0 416 0 1 770
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1681685098
transform 1 0 424 0 1 770
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1681685098
transform 1 0 432 0 1 770
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1681685098
transform 1 0 440 0 1 770
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1681685098
transform 1 0 448 0 1 770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_33
timestamp 1681685098
transform -1 0 512 0 1 770
box -8 -3 64 105
use OR2X1  OR2X1_35
timestamp 1681685098
transform 1 0 512 0 1 770
box -8 -3 40 105
use NOR2X1  NOR2X1_16
timestamp 1681685098
transform 1 0 544 0 1 770
box -8 -3 32 105
use FILL  FILL_1104
timestamp 1681685098
transform 1 0 568 0 1 770
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1681685098
transform 1 0 576 0 1 770
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1681685098
transform 1 0 584 0 1 770
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1681685098
transform 1 0 592 0 1 770
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1681685098
transform 1 0 600 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_17
timestamp 1681685098
transform -1 0 632 0 1 770
box -8 -3 32 105
use FILL  FILL_1115
timestamp 1681685098
transform 1 0 632 0 1 770
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1681685098
transform 1 0 640 0 1 770
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1681685098
transform 1 0 648 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_14
timestamp 1681685098
transform 1 0 656 0 1 770
box -8 -3 40 105
use FILL  FILL_1121
timestamp 1681685098
transform 1 0 688 0 1 770
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1681685098
transform 1 0 696 0 1 770
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1681685098
transform 1 0 704 0 1 770
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1681685098
transform 1 0 712 0 1 770
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1681685098
transform 1 0 720 0 1 770
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1681685098
transform 1 0 728 0 1 770
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1681685098
transform 1 0 736 0 1 770
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1681685098
transform 1 0 744 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_19
timestamp 1681685098
transform -1 0 784 0 1 770
box -8 -3 40 105
use FILL  FILL_1138
timestamp 1681685098
transform 1 0 784 0 1 770
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1681685098
transform 1 0 792 0 1 770
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1681685098
transform 1 0 800 0 1 770
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1681685098
transform 1 0 808 0 1 770
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1681685098
transform 1 0 816 0 1 770
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1681685098
transform 1 0 824 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_5
timestamp 1681685098
transform -1 0 872 0 1 770
box -8 -3 46 105
use FILL  FILL_1145
timestamp 1681685098
transform 1 0 872 0 1 770
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1681685098
transform 1 0 880 0 1 770
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1681685098
transform 1 0 888 0 1 770
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1681685098
transform 1 0 896 0 1 770
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1681685098
transform 1 0 904 0 1 770
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1681685098
transform 1 0 912 0 1 770
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1681685098
transform 1 0 920 0 1 770
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1681685098
transform 1 0 928 0 1 770
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1681685098
transform 1 0 936 0 1 770
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1681685098
transform 1 0 944 0 1 770
box -8 -3 16 105
use INVX2  INVX2_52
timestamp 1681685098
transform 1 0 952 0 1 770
box -9 -3 26 105
use AOI21X1  AOI21X1_6
timestamp 1681685098
transform 1 0 968 0 1 770
box -7 -3 39 105
use FILL  FILL_1166
timestamp 1681685098
transform 1 0 1000 0 1 770
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1681685098
transform 1 0 1008 0 1 770
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1681685098
transform 1 0 1016 0 1 770
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1681685098
transform 1 0 1024 0 1 770
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1681685098
transform 1 0 1032 0 1 770
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1681685098
transform 1 0 1040 0 1 770
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1681685098
transform 1 0 1048 0 1 770
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1681685098
transform 1 0 1056 0 1 770
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1681685098
transform 1 0 1064 0 1 770
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1681685098
transform 1 0 1072 0 1 770
box -8 -3 16 105
use INVX2  INVX2_53
timestamp 1681685098
transform -1 0 1096 0 1 770
box -9 -3 26 105
use AND2X2  AND2X2_22
timestamp 1681685098
transform -1 0 1128 0 1 770
box -8 -3 40 105
use FILL  FILL_1188
timestamp 1681685098
transform 1 0 1128 0 1 770
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1681685098
transform 1 0 1136 0 1 770
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1681685098
transform 1 0 1144 0 1 770
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1681685098
transform 1 0 1152 0 1 770
box -8 -3 16 105
use INVX2  INVX2_54
timestamp 1681685098
transform 1 0 1160 0 1 770
box -9 -3 26 105
use FILL  FILL_1192
timestamp 1681685098
transform 1 0 1176 0 1 770
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1681685098
transform 1 0 1184 0 1 770
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1681685098
transform 1 0 1192 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_23
timestamp 1681685098
transform 1 0 1200 0 1 770
box -8 -3 40 105
use FILL  FILL_1204
timestamp 1681685098
transform 1 0 1232 0 1 770
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1681685098
transform 1 0 1240 0 1 770
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1681685098
transform 1 0 1248 0 1 770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_36
timestamp 1681685098
transform 1 0 1256 0 1 770
box -8 -3 64 105
use OR2X1  OR2X1_37
timestamp 1681685098
transform 1 0 1312 0 1 770
box -8 -3 40 105
use FILL  FILL_1207
timestamp 1681685098
transform 1 0 1344 0 1 770
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1681685098
transform 1 0 1352 0 1 770
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1681685098
transform 1 0 1360 0 1 770
box -8 -3 16 105
use FAX1  FAX1_4
timestamp 1681685098
transform 1 0 1368 0 1 770
box -5 -3 126 105
use FILL  FILL_1210
timestamp 1681685098
transform 1 0 1488 0 1 770
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1681685098
transform 1 0 1496 0 1 770
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1681685098
transform 1 0 1504 0 1 770
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1681685098
transform 1 0 1512 0 1 770
box -8 -3 16 105
use INVX2  INVX2_56
timestamp 1681685098
transform 1 0 1520 0 1 770
box -9 -3 26 105
use FILL  FILL_1214
timestamp 1681685098
transform 1 0 1536 0 1 770
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1681685098
transform 1 0 1544 0 1 770
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1681685098
transform 1 0 1552 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_55
timestamp 1681685098
transform 1 0 1560 0 1 770
box -8 -3 34 105
use FILL  FILL_1243
timestamp 1681685098
transform 1 0 1592 0 1 770
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1681685098
transform 1 0 1600 0 1 770
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1681685098
transform 1 0 1608 0 1 770
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1681685098
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1681685098
transform 1 0 1624 0 1 770
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1681685098
transform 1 0 1632 0 1 770
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1681685098
transform 1 0 1640 0 1 770
box -8 -3 16 105
use BUFX2  BUFX2_12
timestamp 1681685098
transform -1 0 1672 0 1 770
box -5 -3 28 105
use FILL  FILL_1255
timestamp 1681685098
transform 1 0 1672 0 1 770
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1681685098
transform 1 0 1680 0 1 770
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1681685098
transform 1 0 1688 0 1 770
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1681685098
transform 1 0 1696 0 1 770
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1681685098
transform 1 0 1704 0 1 770
box -8 -3 16 105
use BUFX2  BUFX2_13
timestamp 1681685098
transform 1 0 1712 0 1 770
box -5 -3 28 105
use FILL  FILL_1265
timestamp 1681685098
transform 1 0 1736 0 1 770
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1681685098
transform 1 0 1744 0 1 770
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1681685098
transform 1 0 1752 0 1 770
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1681685098
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1681685098
transform 1 0 1768 0 1 770
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1681685098
transform 1 0 1776 0 1 770
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1681685098
transform 1 0 1784 0 1 770
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1681685098
transform 1 0 1792 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_42
timestamp 1681685098
transform 1 0 1800 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1681685098
transform -1 0 1848 0 1 770
box -8 -3 32 105
use FILL  FILL_1280
timestamp 1681685098
transform 1 0 1848 0 1 770
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1681685098
transform 1 0 1856 0 1 770
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1681685098
transform 1 0 1864 0 1 770
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1681685098
transform 1 0 1872 0 1 770
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1681685098
transform 1 0 1880 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1681685098
transform 1 0 1888 0 1 770
box -8 -3 104 105
use FILL  FILL_1288
timestamp 1681685098
transform 1 0 1984 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_20
timestamp 1681685098
transform 1 0 1992 0 1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_56
timestamp 1681685098
transform 1 0 2016 0 1 770
box -8 -3 34 105
use FILL  FILL_1289
timestamp 1681685098
transform 1 0 2048 0 1 770
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1681685098
transform 1 0 2056 0 1 770
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1681685098
transform 1 0 2064 0 1 770
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1681685098
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1681685098
transform 1 0 2080 0 1 770
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1681685098
transform 1 0 2088 0 1 770
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1681685098
transform 1 0 2096 0 1 770
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1681685098
transform 1 0 2104 0 1 770
box -8 -3 16 105
use INVX2  INVX2_59
timestamp 1681685098
transform -1 0 2128 0 1 770
box -9 -3 26 105
use FILL  FILL_1297
timestamp 1681685098
transform 1 0 2128 0 1 770
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1681685098
transform 1 0 2136 0 1 770
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_25
timestamp 1681685098
transform 1 0 2170 0 1 770
box -10 -3 10 3
use M3_M2  M3_M2_746
timestamp 1681685098
transform 1 0 100 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1681685098
transform 1 0 132 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1681685098
transform 1 0 124 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1092
timestamp 1681685098
transform 1 0 84 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1681685098
transform 1 0 132 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_754
timestamp 1681685098
transform 1 0 156 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1681685098
transform 1 0 172 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1094
timestamp 1681685098
transform 1 0 180 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1681685098
transform 1 0 148 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1681685098
transform 1 0 156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1681685098
transform 1 0 172 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_789
timestamp 1681685098
transform 1 0 148 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1681685098
transform 1 0 172 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1681685098
transform 1 0 236 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1095
timestamp 1681685098
transform 1 0 236 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_764
timestamp 1681685098
transform 1 0 268 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1135
timestamp 1681685098
transform 1 0 260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1681685098
transform 1 0 276 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_755
timestamp 1681685098
transform 1 0 372 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1681685098
transform 1 0 300 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1681685098
transform 1 0 364 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1681685098
transform 1 0 404 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1097
timestamp 1681685098
transform 1 0 388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1681685098
transform 1 0 404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1681685098
transform 1 0 284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1681685098
transform 1 0 300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1681685098
transform 1 0 308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1681685098
transform 1 0 364 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_791
timestamp 1681685098
transform 1 0 284 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1681685098
transform 1 0 308 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1173
timestamp 1681685098
transform 1 0 404 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1681685098
transform 1 0 428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1681685098
transform 1 0 444 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_780
timestamp 1681685098
transform 1 0 444 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1681685098
transform 1 0 436 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1681685098
transform 1 0 476 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1681685098
transform 1 0 548 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_1086
timestamp 1681685098
transform 1 0 476 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_768
timestamp 1681685098
transform 1 0 484 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1681685098
transform 1 0 508 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1101
timestamp 1681685098
transform 1 0 484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1681685098
transform 1 0 508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1681685098
transform 1 0 500 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_781
timestamp 1681685098
transform 1 0 508 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1681685098
transform 1 0 556 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1103
timestamp 1681685098
transform 1 0 556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1681685098
transform 1 0 564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1681685098
transform 1 0 540 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_794
timestamp 1681685098
transform 1 0 540 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1105
timestamp 1681685098
transform 1 0 628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1681685098
transform 1 0 612 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_782
timestamp 1681685098
transform 1 0 628 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1681685098
transform 1 0 612 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1681685098
transform 1 0 660 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_1087
timestamp 1681685098
transform 1 0 652 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1681685098
transform 1 0 644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1681685098
transform 1 0 780 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_778
timestamp 1681685098
transform 1 0 788 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1108
timestamp 1681685098
transform 1 0 812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1681685098
transform 1 0 748 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1681685098
transform 1 0 756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1681685098
transform 1 0 772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1681685098
transform 1 0 788 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1681685098
transform 1 0 804 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_795
timestamp 1681685098
transform 1 0 748 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1681685098
transform 1 0 772 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1681685098
transform 1 0 812 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1681685098
transform 1 0 804 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1681685098
transform 1 0 852 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1109
timestamp 1681685098
transform 1 0 852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1681685098
transform 1 0 844 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1681685098
transform 1 0 860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1681685098
transform 1 0 876 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_796
timestamp 1681685098
transform 1 0 860 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1681685098
transform 1 0 972 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1681685098
transform 1 0 964 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1088
timestamp 1681685098
transform 1 0 972 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1681685098
transform 1 0 972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1681685098
transform 1 0 988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1681685098
transform 1 0 964 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1681685098
transform 1 0 1004 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_759
timestamp 1681685098
transform 1 0 1100 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1681685098
transform 1 0 1092 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1112
timestamp 1681685098
transform 1 0 1092 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1681685098
transform 1 0 1100 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_821
timestamp 1681685098
transform 1 0 1116 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_1174
timestamp 1681685098
transform 1 0 1140 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1681685098
transform 1 0 1180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1681685098
transform 1 0 1220 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1681685098
transform 1 0 1220 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_797
timestamp 1681685098
transform 1 0 1220 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1154
timestamp 1681685098
transform 1 0 1244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1681685098
transform 1 0 1260 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_798
timestamp 1681685098
transform 1 0 1260 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1681685098
transform 1 0 1244 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1681685098
transform 1 0 1364 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1115
timestamp 1681685098
transform 1 0 1364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1681685098
transform 1 0 1340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1681685098
transform 1 0 1348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1681685098
transform 1 0 1364 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_811
timestamp 1681685098
transform 1 0 1364 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_1184
timestamp 1681685098
transform 1 0 1372 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1681685098
transform 1 0 1396 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_812
timestamp 1681685098
transform 1 0 1396 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1681685098
transform 1 0 1420 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1176
timestamp 1681685098
transform 1 0 1420 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1681685098
transform 1 0 1436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1681685098
transform 1 0 1444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1681685098
transform 1 0 1436 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1681685098
transform 1 0 1492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1681685098
transform 1 0 1492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1681685098
transform 1 0 1516 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_799
timestamp 1681685098
transform 1 0 1484 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1178
timestamp 1681685098
transform 1 0 1500 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_800
timestamp 1681685098
transform 1 0 1508 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1179
timestamp 1681685098
transform 1 0 1516 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_813
timestamp 1681685098
transform 1 0 1500 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_1185
timestamp 1681685098
transform 1 0 1508 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1681685098
transform 1 0 1532 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_784
timestamp 1681685098
transform 1 0 1532 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1120
timestamp 1681685098
transform 1 0 1620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1681685098
transform 1 0 1628 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_801
timestamp 1681685098
transform 1 0 1628 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1180
timestamp 1681685098
transform 1 0 1644 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_822
timestamp 1681685098
transform 1 0 1644 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_1121
timestamp 1681685098
transform 1 0 1668 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_774
timestamp 1681685098
transform 1 0 1684 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1162
timestamp 1681685098
transform 1 0 1684 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_750
timestamp 1681685098
transform 1 0 1708 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1681685098
transform 1 0 1700 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_1122
timestamp 1681685098
transform 1 0 1716 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1681685098
transform 1 0 1708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1681685098
transform 1 0 1708 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_819
timestamp 1681685098
transform 1 0 1692 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_1090
timestamp 1681685098
transform 1 0 1740 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1681685098
transform 1 0 1732 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_802
timestamp 1681685098
transform 1 0 1732 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1681685098
transform 1 0 1740 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_1091
timestamp 1681685098
transform 1 0 1756 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1681685098
transform 1 0 1812 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_803
timestamp 1681685098
transform 1 0 1820 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1681685098
transform 1 0 1836 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1124
timestamp 1681685098
transform 1 0 1828 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1681685098
transform 1 0 1836 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_785
timestamp 1681685098
transform 1 0 1828 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1681685098
transform 1 0 1844 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1126
timestamp 1681685098
transform 1 0 1852 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_786
timestamp 1681685098
transform 1 0 1852 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1681685098
transform 1 0 1868 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1165
timestamp 1681685098
transform 1 0 1860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1681685098
transform 1 0 1868 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_814
timestamp 1681685098
transform 1 0 1860 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1681685098
transform 1 0 1924 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_1127
timestamp 1681685098
transform 1 0 1900 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1681685098
transform 1 0 1908 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_787
timestamp 1681685098
transform 1 0 1900 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1182
timestamp 1681685098
transform 1 0 1900 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1681685098
transform 1 0 2004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1681685098
transform 1 0 1916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1681685098
transform 1 0 1924 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_788
timestamp 1681685098
transform 1 0 1940 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_1169
timestamp 1681685098
transform 1 0 1956 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_804
timestamp 1681685098
transform 1 0 1916 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1681685098
transform 1 0 1956 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1681685098
transform 1 0 2028 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1681685098
transform 1 0 2108 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_1130
timestamp 1681685098
transform 1 0 2028 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_777
timestamp 1681685098
transform 1 0 2132 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_1131
timestamp 1681685098
transform 1 0 2132 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1681685098
transform 1 0 2052 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1681685098
transform 1 0 2116 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1681685098
transform 1 0 2124 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_806
timestamp 1681685098
transform 1 0 2068 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_1183
timestamp 1681685098
transform 1 0 2116 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_807
timestamp 1681685098
transform 1 0 2124 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1681685098
transform 1 0 2108 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1681685098
transform 1 0 2124 0 1 705
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_26
timestamp 1681685098
transform 1 0 24 0 1 670
box -10 -3 10 3
use FILL  FILL_1078
timestamp 1681685098
transform 1 0 72 0 -1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_11
timestamp 1681685098
transform 1 0 80 0 -1 770
box -8 -3 64 105
use FILL  FILL_1083
timestamp 1681685098
transform 1 0 136 0 -1 770
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1681685098
transform 1 0 144 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_17
timestamp 1681685098
transform -1 0 184 0 -1 770
box -8 -3 40 105
use XOR2X1  XOR2X1_13
timestamp 1681685098
transform 1 0 184 0 -1 770
box -8 -3 64 105
use FILL  FILL_1087
timestamp 1681685098
transform 1 0 240 0 -1 770
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1681685098
transform 1 0 248 0 -1 770
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1681685098
transform 1 0 256 0 -1 770
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1681685098
transform 1 0 264 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_18
timestamp 1681685098
transform 1 0 272 0 -1 770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1681685098
transform -1 0 400 0 -1 770
box -8 -3 104 105
use OAI21X1  OAI21X1_51
timestamp 1681685098
transform -1 0 432 0 -1 770
box -8 -3 34 105
use INVX2  INVX2_51
timestamp 1681685098
transform -1 0 448 0 -1 770
box -9 -3 26 105
use FILL  FILL_1106
timestamp 1681685098
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1681685098
transform 1 0 456 0 -1 770
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1681685098
transform 1 0 464 0 -1 770
box -8 -3 16 105
use OR2X1  OR2X1_36
timestamp 1681685098
transform 1 0 472 0 -1 770
box -8 -3 40 105
use XNOR2X1  XNOR2X1_34
timestamp 1681685098
transform 1 0 504 0 -1 770
box -8 -3 64 105
use FILL  FILL_1109
timestamp 1681685098
transform 1 0 560 0 -1 770
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1681685098
transform 1 0 568 0 -1 770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_35
timestamp 1681685098
transform 1 0 576 0 -1 770
box -8 -3 64 105
use FILL  FILL_1116
timestamp 1681685098
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1681685098
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1681685098
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1681685098
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1681685098
transform 1 0 664 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_18
timestamp 1681685098
transform 1 0 672 0 -1 770
box -8 -3 32 105
use FILL  FILL_1125
timestamp 1681685098
transform 1 0 696 0 -1 770
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1681685098
transform 1 0 704 0 -1 770
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1681685098
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1681685098
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1681685098
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1681685098
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1681685098
transform 1 0 744 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_20
timestamp 1681685098
transform -1 0 784 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1681685098
transform -1 0 816 0 -1 770
box -8 -3 40 105
use FILL  FILL_1143
timestamp 1681685098
transform 1 0 816 0 -1 770
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1681685098
transform 1 0 824 0 -1 770
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1681685098
transform 1 0 832 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_6
timestamp 1681685098
transform 1 0 840 0 -1 770
box -8 -3 46 105
use FILL  FILL_1149
timestamp 1681685098
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1681685098
transform 1 0 888 0 -1 770
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1681685098
transform 1 0 896 0 -1 770
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1681685098
transform 1 0 904 0 -1 770
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1681685098
transform 1 0 912 0 -1 770
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1681685098
transform 1 0 920 0 -1 770
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1681685098
transform 1 0 928 0 -1 770
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1681685098
transform 1 0 936 0 -1 770
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1681685098
transform 1 0 944 0 -1 770
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1681685098
transform 1 0 952 0 -1 770
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1681685098
transform 1 0 960 0 -1 770
box -8 -3 16 105
use AOI21X1  AOI21X1_7
timestamp 1681685098
transform -1 0 1000 0 -1 770
box -7 -3 39 105
use FILL  FILL_1169
timestamp 1681685098
transform 1 0 1000 0 -1 770
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1681685098
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1681685098
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1681685098
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1681685098
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1681685098
transform 1 0 1040 0 -1 770
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1681685098
transform 1 0 1048 0 -1 770
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1681685098
transform 1 0 1056 0 -1 770
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1681685098
transform 1 0 1064 0 -1 770
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1681685098
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_55
timestamp 1681685098
transform -1 0 1096 0 -1 770
box -9 -3 26 105
use FILL  FILL_1193
timestamp 1681685098
transform 1 0 1096 0 -1 770
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1681685098
transform 1 0 1104 0 -1 770
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1681685098
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1681685098
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1681685098
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_52
timestamp 1681685098
transform -1 0 1168 0 -1 770
box -8 -3 34 105
use FILL  FILL_1198
timestamp 1681685098
transform 1 0 1168 0 -1 770
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1681685098
transform 1 0 1176 0 -1 770
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1681685098
transform 1 0 1184 0 -1 770
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1681685098
transform 1 0 1192 0 -1 770
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1681685098
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1681685098
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1681685098
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1681685098
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_24
timestamp 1681685098
transform 1 0 1232 0 -1 770
box -8 -3 40 105
use FILL  FILL_1219
timestamp 1681685098
transform 1 0 1264 0 -1 770
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1681685098
transform 1 0 1272 0 -1 770
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1681685098
transform 1 0 1280 0 -1 770
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1681685098
transform 1 0 1288 0 -1 770
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1681685098
transform 1 0 1296 0 -1 770
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1681685098
transform 1 0 1304 0 -1 770
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1681685098
transform 1 0 1312 0 -1 770
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1681685098
transform 1 0 1320 0 -1 770
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1681685098
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_823
timestamp 1681685098
transform 1 0 1364 0 1 675
box -3 -3 3 3
use OAI21X1  OAI21X1_53
timestamp 1681685098
transform 1 0 1336 0 -1 770
box -8 -3 34 105
use FILL  FILL_1228
timestamp 1681685098
transform 1 0 1368 0 -1 770
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1681685098
transform 1 0 1376 0 -1 770
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1681685098
transform 1 0 1384 0 -1 770
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1681685098
transform 1 0 1392 0 -1 770
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1681685098
transform 1 0 1400 0 -1 770
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1681685098
transform 1 0 1408 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_824
timestamp 1681685098
transform 1 0 1436 0 1 675
box -3 -3 3 3
use NAND2X1  NAND2X1_39
timestamp 1681685098
transform -1 0 1440 0 -1 770
box -8 -3 32 105
use FILL  FILL_1234
timestamp 1681685098
transform 1 0 1440 0 -1 770
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1681685098
transform 1 0 1448 0 -1 770
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1681685098
transform 1 0 1456 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_54
timestamp 1681685098
transform -1 0 1496 0 -1 770
box -8 -3 34 105
use M3_M2  M3_M2_825
timestamp 1681685098
transform 1 0 1516 0 1 675
box -3 -3 3 3
use NAND3X1  NAND3X1_15
timestamp 1681685098
transform -1 0 1528 0 -1 770
box -8 -3 40 105
use FILL  FILL_1237
timestamp 1681685098
transform 1 0 1528 0 -1 770
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1681685098
transform 1 0 1536 0 -1 770
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1681685098
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1681685098
transform 1 0 1552 0 -1 770
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1681685098
transform 1 0 1560 0 -1 770
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1681685098
transform 1 0 1568 0 -1 770
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1681685098
transform 1 0 1576 0 -1 770
box -8 -3 16 105
use BUFX2  BUFX2_11
timestamp 1681685098
transform -1 0 1608 0 -1 770
box -5 -3 28 105
use FILL  FILL_1249
timestamp 1681685098
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1681685098
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_40
timestamp 1681685098
transform 1 0 1624 0 -1 770
box -8 -3 32 105
use FILL  FILL_1256
timestamp 1681685098
transform 1 0 1648 0 -1 770
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1681685098
transform 1 0 1656 0 -1 770
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1681685098
transform 1 0 1664 0 -1 770
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1681685098
transform 1 0 1672 0 -1 770
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1681685098
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_41
timestamp 1681685098
transform 1 0 1688 0 -1 770
box -8 -3 32 105
use BUFX2  BUFX2_14
timestamp 1681685098
transform -1 0 1736 0 -1 770
box -5 -3 28 105
use FILL  FILL_1266
timestamp 1681685098
transform 1 0 1736 0 -1 770
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1681685098
transform 1 0 1744 0 -1 770
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1681685098
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1681685098
transform 1 0 1760 0 -1 770
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1681685098
transform 1 0 1768 0 -1 770
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1681685098
transform 1 0 1776 0 -1 770
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1681685098
transform 1 0 1784 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_19
timestamp 1681685098
transform 1 0 1792 0 -1 770
box -8 -3 32 105
use INVX2  INVX2_57
timestamp 1681685098
transform -1 0 1832 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1681685098
transform 1 0 1832 0 -1 770
box -9 -3 26 105
use FILL  FILL_1281
timestamp 1681685098
transform 1 0 1848 0 -1 770
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1681685098
transform 1 0 1856 0 -1 770
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1681685098
transform 1 0 1864 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_57
timestamp 1681685098
transform 1 0 1872 0 -1 770
box -8 -3 34 105
use INVX2  INVX2_60
timestamp 1681685098
transform 1 0 1904 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1681685098
transform -1 0 2016 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1681685098
transform 1 0 2016 0 -1 770
box -8 -3 104 105
use NAND2X1  NAND2X1_44
timestamp 1681685098
transform -1 0 2136 0 -1 770
box -8 -3 32 105
use FILL  FILL_1299
timestamp 1681685098
transform 1 0 2136 0 -1 770
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_27
timestamp 1681685098
transform 1 0 2194 0 1 670
box -10 -3 10 3
use M2_M1  M2_M1_1191
timestamp 1681685098
transform 1 0 84 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_859
timestamp 1681685098
transform 1 0 84 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_1192
timestamp 1681685098
transform 1 0 108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1681685098
transform 1 0 116 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_860
timestamp 1681685098
transform 1 0 116 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1681685098
transform 1 0 132 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1681685098
transform 1 0 156 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1681685098
transform 1 0 180 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1681685098
transform 1 0 212 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1193
timestamp 1681685098
transform 1 0 156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1681685098
transform 1 0 172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1681685098
transform 1 0 188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1681685098
transform 1 0 212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1681685098
transform 1 0 180 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_861
timestamp 1681685098
transform 1 0 180 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1681685098
transform 1 0 300 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_1197
timestamp 1681685098
transform 1 0 252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1681685098
transform 1 0 276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1681685098
transform 1 0 300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1681685098
transform 1 0 308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1681685098
transform 1 0 236 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1681685098
transform 1 0 244 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_862
timestamp 1681685098
transform 1 0 236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1681685098
transform 1 0 268 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_1235
timestamp 1681685098
transform 1 0 332 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_864
timestamp 1681685098
transform 1 0 332 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1681685098
transform 1 0 380 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1681685098
transform 1 0 404 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1201
timestamp 1681685098
transform 1 0 372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1681685098
transform 1 0 380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1681685098
transform 1 0 396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1681685098
transform 1 0 412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1681685098
transform 1 0 388 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_869
timestamp 1681685098
transform 1 0 388 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1681685098
transform 1 0 404 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1681685098
transform 1 0 428 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1205
timestamp 1681685098
transform 1 0 428 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_850
timestamp 1681685098
transform 1 0 444 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1681685098
transform 1 0 452 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1681685098
transform 1 0 468 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_1237
timestamp 1681685098
transform 1 0 468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1681685098
transform 1 0 484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1681685098
transform 1 0 508 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_843
timestamp 1681685098
transform 1 0 532 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1238
timestamp 1681685098
transform 1 0 532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1681685098
transform 1 0 532 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_872
timestamp 1681685098
transform 1 0 532 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1681685098
transform 1 0 612 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1681685098
transform 1 0 564 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1207
timestamp 1681685098
transform 1 0 564 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_851
timestamp 1681685098
transform 1 0 596 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1208
timestamp 1681685098
transform 1 0 604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1681685098
transform 1 0 548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1681685098
transform 1 0 572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1681685098
transform 1 0 620 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_865
timestamp 1681685098
transform 1 0 620 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_1242
timestamp 1681685098
transform 1 0 636 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_828
timestamp 1681685098
transform 1 0 700 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_1209
timestamp 1681685098
transform 1 0 676 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_852
timestamp 1681685098
transform 1 0 684 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1210
timestamp 1681685098
transform 1 0 692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1681685098
transform 1 0 700 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_832
timestamp 1681685098
transform 1 0 740 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_1244
timestamp 1681685098
transform 1 0 764 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_833
timestamp 1681685098
transform 1 0 788 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_1186
timestamp 1681685098
transform 1 0 812 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_845
timestamp 1681685098
transform 1 0 844 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1211
timestamp 1681685098
transform 1 0 860 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_873
timestamp 1681685098
transform 1 0 860 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_1212
timestamp 1681685098
transform 1 0 876 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_846
timestamp 1681685098
transform 1 0 892 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1213
timestamp 1681685098
transform 1 0 892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1681685098
transform 1 0 884 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_834
timestamp 1681685098
transform 1 0 964 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_1246
timestamp 1681685098
transform 1 0 964 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1681685098
transform 1 0 972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1681685098
transform 1 0 988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1681685098
transform 1 0 1052 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_829
timestamp 1681685098
transform 1 0 1116 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1681685098
transform 1 0 1132 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1248
timestamp 1681685098
transform 1 0 1132 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1681685098
transform 1 0 1140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1681685098
transform 1 0 1156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1681685098
transform 1 0 1180 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1681685098
transform 1 0 1220 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_848
timestamp 1681685098
transform 1 0 1252 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1216
timestamp 1681685098
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1681685098
transform 1 0 1332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1681685098
transform 1 0 1348 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1681685098
transform 1 0 1348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1681685098
transform 1 0 1364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1681685098
transform 1 0 1388 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_835
timestamp 1681685098
transform 1 0 1444 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_1218
timestamp 1681685098
transform 1 0 1412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1681685098
transform 1 0 1508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1681685098
transform 1 0 1516 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_866
timestamp 1681685098
transform 1 0 1404 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_1259
timestamp 1681685098
transform 1 0 1500 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_867
timestamp 1681685098
transform 1 0 1508 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_1256
timestamp 1681685098
transform 1 0 1628 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1681685098
transform 1 0 1676 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1681685098
transform 1 0 1764 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_857
timestamp 1681685098
transform 1 0 1764 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1681685098
transform 1 0 1780 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1220
timestamp 1681685098
transform 1 0 1804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1681685098
transform 1 0 1860 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1681685098
transform 1 0 1780 0 1 607
box -2 -2 2 2
use M3_M2  M3_M2_868
timestamp 1681685098
transform 1 0 1860 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1681685098
transform 1 0 1996 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1681685098
transform 1 0 1916 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1222
timestamp 1681685098
transform 1 0 1940 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_855
timestamp 1681685098
transform 1 0 1988 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_1223
timestamp 1681685098
transform 1 0 1996 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1681685098
transform 1 0 1916 0 1 607
box -2 -2 2 2
use M3_M2  M3_M2_858
timestamp 1681685098
transform 1 0 1956 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1681685098
transform 1 0 2036 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1681685098
transform 1 0 2148 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_1224
timestamp 1681685098
transform 1 0 2060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1681685098
transform 1 0 2116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1681685098
transform 1 0 2124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1681685098
transform 1 0 2036 0 1 607
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1681685098
transform 1 0 2148 0 1 615
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_28
timestamp 1681685098
transform 1 0 48 0 1 570
box -10 -3 10 3
use FILL  FILL_1300
timestamp 1681685098
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1681685098
transform 1 0 80 0 1 570
box -8 -3 16 105
use AND2X2  AND2X2_25
timestamp 1681685098
transform -1 0 120 0 1 570
box -8 -3 40 105
use FILL  FILL_1303
timestamp 1681685098
transform 1 0 120 0 1 570
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1681685098
transform 1 0 128 0 1 570
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1681685098
transform 1 0 136 0 1 570
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1681685098
transform 1 0 144 0 1 570
box -8 -3 16 105
use AND2X2  AND2X2_26
timestamp 1681685098
transform -1 0 184 0 1 570
box -8 -3 40 105
use XOR2X1  XOR2X1_15
timestamp 1681685098
transform -1 0 240 0 1 570
box -8 -3 64 105
use AND2X2  AND2X2_27
timestamp 1681685098
transform 1 0 240 0 1 570
box -8 -3 40 105
use XOR2X1  XOR2X1_16
timestamp 1681685098
transform 1 0 272 0 1 570
box -8 -3 64 105
use FILL  FILL_1315
timestamp 1681685098
transform 1 0 328 0 1 570
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1681685098
transform 1 0 336 0 1 570
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1681685098
transform 1 0 344 0 1 570
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1681685098
transform 1 0 352 0 1 570
box -8 -3 16 105
use INVX2  INVX2_61
timestamp 1681685098
transform 1 0 360 0 1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_7
timestamp 1681685098
transform -1 0 416 0 1 570
box -8 -3 46 105
use FILL  FILL_1319
timestamp 1681685098
transform 1 0 416 0 1 570
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1681685098
transform 1 0 424 0 1 570
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1681685098
transform 1 0 432 0 1 570
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1681685098
transform 1 0 440 0 1 570
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1681685098
transform 1 0 448 0 1 570
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1681685098
transform 1 0 456 0 1 570
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1681685098
transform 1 0 464 0 1 570
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1681685098
transform 1 0 472 0 1 570
box -8 -3 16 105
use OR2X1  OR2X1_38
timestamp 1681685098
transform -1 0 512 0 1 570
box -8 -3 40 105
use FILL  FILL_1333
timestamp 1681685098
transform 1 0 512 0 1 570
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1681685098
transform 1 0 520 0 1 570
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1681685098
transform 1 0 528 0 1 570
box -8 -3 16 105
use OR2X1  OR2X1_39
timestamp 1681685098
transform 1 0 536 0 1 570
box -8 -3 40 105
use XNOR2X1  XNOR2X1_37
timestamp 1681685098
transform 1 0 568 0 1 570
box -8 -3 64 105
use FILL  FILL_1336
timestamp 1681685098
transform 1 0 624 0 1 570
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1681685098
transform 1 0 632 0 1 570
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1681685098
transform 1 0 640 0 1 570
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1681685098
transform 1 0 648 0 1 570
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1681685098
transform 1 0 656 0 1 570
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1681685098
transform 1 0 664 0 1 570
box -8 -3 16 105
use AND2X2  AND2X2_29
timestamp 1681685098
transform -1 0 704 0 1 570
box -8 -3 40 105
use FILL  FILL_1346
timestamp 1681685098
transform 1 0 704 0 1 570
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1681685098
transform 1 0 712 0 1 570
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1681685098
transform 1 0 720 0 1 570
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1681685098
transform 1 0 728 0 1 570
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1681685098
transform 1 0 736 0 1 570
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1681685098
transform 1 0 744 0 1 570
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1681685098
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1681685098
transform 1 0 760 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_45
timestamp 1681685098
transform 1 0 768 0 1 570
box -8 -3 32 105
use FILL  FILL_1354
timestamp 1681685098
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1681685098
transform 1 0 800 0 1 570
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1681685098
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1681685098
transform 1 0 816 0 1 570
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1681685098
transform 1 0 824 0 1 570
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1681685098
transform 1 0 832 0 1 570
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1681685098
transform 1 0 840 0 1 570
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1681685098
transform 1 0 848 0 1 570
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1681685098
transform 1 0 856 0 1 570
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1681685098
transform 1 0 864 0 1 570
box -8 -3 16 105
use INVX2  INVX2_62
timestamp 1681685098
transform -1 0 888 0 1 570
box -9 -3 26 105
use FILL  FILL_1371
timestamp 1681685098
transform 1 0 888 0 1 570
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1681685098
transform 1 0 896 0 1 570
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1681685098
transform 1 0 904 0 1 570
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1681685098
transform 1 0 912 0 1 570
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1681685098
transform 1 0 920 0 1 570
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1681685098
transform 1 0 928 0 1 570
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1681685098
transform 1 0 936 0 1 570
box -8 -3 16 105
use AOI21X1  AOI21X1_8
timestamp 1681685098
transform -1 0 976 0 1 570
box -7 -3 39 105
use FILL  FILL_1382
timestamp 1681685098
transform 1 0 976 0 1 570
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1681685098
transform 1 0 984 0 1 570
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1681685098
transform 1 0 992 0 1 570
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1681685098
transform 1 0 1000 0 1 570
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1681685098
transform 1 0 1008 0 1 570
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1681685098
transform 1 0 1016 0 1 570
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1681685098
transform 1 0 1024 0 1 570
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1681685098
transform 1 0 1032 0 1 570
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1681685098
transform 1 0 1040 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_59
timestamp 1681685098
transform -1 0 1080 0 1 570
box -8 -3 34 105
use FILL  FILL_1391
timestamp 1681685098
transform 1 0 1080 0 1 570
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1681685098
transform 1 0 1088 0 1 570
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1681685098
transform 1 0 1096 0 1 570
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1681685098
transform 1 0 1104 0 1 570
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1681685098
transform 1 0 1112 0 1 570
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1681685098
transform 1 0 1120 0 1 570
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1681685098
transform 1 0 1128 0 1 570
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1681685098
transform 1 0 1136 0 1 570
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1681685098
transform 1 0 1144 0 1 570
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1681685098
transform 1 0 1152 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_48
timestamp 1681685098
transform 1 0 1160 0 1 570
box -8 -3 32 105
use FILL  FILL_1412
timestamp 1681685098
transform 1 0 1184 0 1 570
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1681685098
transform 1 0 1192 0 1 570
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1681685098
transform 1 0 1200 0 1 570
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1681685098
transform 1 0 1208 0 1 570
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1681685098
transform 1 0 1216 0 1 570
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1681685098
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1681685098
transform 1 0 1232 0 1 570
box -8 -3 16 105
use INVX2  INVX2_63
timestamp 1681685098
transform 1 0 1240 0 1 570
box -9 -3 26 105
use FILL  FILL_1425
timestamp 1681685098
transform 1 0 1256 0 1 570
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1681685098
transform 1 0 1264 0 1 570
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1681685098
transform 1 0 1272 0 1 570
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1681685098
transform 1 0 1280 0 1 570
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1681685098
transform 1 0 1288 0 1 570
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1681685098
transform 1 0 1296 0 1 570
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1681685098
transform 1 0 1304 0 1 570
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1681685098
transform 1 0 1312 0 1 570
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1681685098
transform 1 0 1320 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_50
timestamp 1681685098
transform 1 0 1328 0 1 570
box -8 -3 32 105
use FILL  FILL_1439
timestamp 1681685098
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1681685098
transform 1 0 1360 0 1 570
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1681685098
transform 1 0 1368 0 1 570
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1681685098
transform 1 0 1376 0 1 570
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1681685098
transform 1 0 1384 0 1 570
box -8 -3 16 105
use FAX1  FAX1_5
timestamp 1681685098
transform 1 0 1392 0 1 570
box -5 -3 126 105
use FILL  FILL_1444
timestamp 1681685098
transform 1 0 1512 0 1 570
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1681685098
transform 1 0 1520 0 1 570
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1681685098
transform 1 0 1528 0 1 570
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1681685098
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1681685098
transform 1 0 1544 0 1 570
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1681685098
transform 1 0 1552 0 1 570
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1681685098
transform 1 0 1560 0 1 570
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1681685098
transform 1 0 1568 0 1 570
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1681685098
transform 1 0 1576 0 1 570
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1681685098
transform 1 0 1584 0 1 570
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1681685098
transform 1 0 1592 0 1 570
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1681685098
transform 1 0 1600 0 1 570
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1681685098
transform 1 0 1608 0 1 570
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1681685098
transform 1 0 1616 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_51
timestamp 1681685098
transform 1 0 1624 0 1 570
box -8 -3 32 105
use FILL  FILL_1466
timestamp 1681685098
transform 1 0 1648 0 1 570
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1681685098
transform 1 0 1656 0 1 570
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1681685098
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1681685098
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1681685098
transform 1 0 1680 0 1 570
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1681685098
transform 1 0 1688 0 1 570
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1681685098
transform 1 0 1696 0 1 570
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1681685098
transform 1 0 1704 0 1 570
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1681685098
transform 1 0 1712 0 1 570
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1681685098
transform 1 0 1720 0 1 570
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1681685098
transform 1 0 1728 0 1 570
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1681685098
transform 1 0 1736 0 1 570
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1681685098
transform 1 0 1744 0 1 570
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1681685098
transform 1 0 1752 0 1 570
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1681685098
transform 1 0 1760 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1681685098
transform 1 0 1768 0 1 570
box -8 -3 104 105
use FILL  FILL_1492
timestamp 1681685098
transform 1 0 1864 0 1 570
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1681685098
transform 1 0 1872 0 1 570
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1681685098
transform 1 0 1880 0 1 570
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1681685098
transform 1 0 1888 0 1 570
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1681685098
transform 1 0 1896 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1681685098
transform 1 0 1904 0 1 570
box -8 -3 104 105
use FILL  FILL_1508
timestamp 1681685098
transform 1 0 2000 0 1 570
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1681685098
transform 1 0 2008 0 1 570
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1681685098
transform 1 0 2016 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_874
timestamp 1681685098
transform 1 0 2036 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1681685098
transform 1 0 2116 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_61
timestamp 1681685098
transform 1 0 2024 0 1 570
box -8 -3 104 105
use INVX2  INVX2_67
timestamp 1681685098
transform 1 0 2120 0 1 570
box -9 -3 26 105
use FILL  FILL_1511
timestamp 1681685098
transform 1 0 2136 0 1 570
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_29
timestamp 1681685098
transform 1 0 2170 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_926
timestamp 1681685098
transform 1 0 108 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1681685098
transform 1 0 132 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1264
timestamp 1681685098
transform 1 0 172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1681685098
transform 1 0 196 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_914
timestamp 1681685098
transform 1 0 172 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1681685098
transform 1 0 196 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1265
timestamp 1681685098
transform 1 0 228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1681685098
transform 1 0 236 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_929
timestamp 1681685098
transform 1 0 228 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1681685098
transform 1 0 324 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1681685098
transform 1 0 364 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1267
timestamp 1681685098
transform 1 0 348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1681685098
transform 1 0 364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1681685098
transform 1 0 244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1681685098
transform 1 0 260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1681685098
transform 1 0 268 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1681685098
transform 1 0 324 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_900
timestamp 1681685098
transform 1 0 348 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1681685098
transform 1 0 260 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1681685098
transform 1 0 268 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1681685098
transform 1 0 244 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1681685098
transform 1 0 268 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_1269
timestamp 1681685098
transform 1 0 396 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1681685098
transform 1 0 404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1681685098
transform 1 0 380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1681685098
transform 1 0 388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1681685098
transform 1 0 412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1681685098
transform 1 0 428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1681685098
transform 1 0 364 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_931
timestamp 1681685098
transform 1 0 364 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1681685098
transform 1 0 412 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1681685098
transform 1 0 412 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_1271
timestamp 1681685098
transform 1 0 444 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_878
timestamp 1681685098
transform 1 0 460 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1272
timestamp 1681685098
transform 1 0 460 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_901
timestamp 1681685098
transform 1 0 460 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1681685098
transform 1 0 564 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1260
timestamp 1681685098
transform 1 0 572 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1681685098
transform 1 0 484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1681685098
transform 1 0 540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1681685098
transform 1 0 548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1681685098
transform 1 0 580 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_944
timestamp 1681685098
transform 1 0 564 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1681685098
transform 1 0 628 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1274
timestamp 1681685098
transform 1 0 628 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_902
timestamp 1681685098
transform 1 0 604 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1309
timestamp 1681685098
transform 1 0 612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1681685098
transform 1 0 628 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_916
timestamp 1681685098
transform 1 0 612 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1681685098
transform 1 0 652 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1681685098
transform 1 0 660 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1681685098
transform 1 0 692 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1261
timestamp 1681685098
transform 1 0 708 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1681685098
transform 1 0 692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1681685098
transform 1 0 716 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_904
timestamp 1681685098
transform 1 0 716 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1681685098
transform 1 0 812 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1276
timestamp 1681685098
transform 1 0 812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1681685098
transform 1 0 732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1681685098
transform 1 0 788 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1681685098
transform 1 0 700 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_917
timestamp 1681685098
transform 1 0 764 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1681685098
transform 1 0 828 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1345
timestamp 1681685098
transform 1 0 828 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1681685098
transform 1 0 884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1681685098
transform 1 0 916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1681685098
transform 1 0 932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1681685098
transform 1 0 948 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_880
timestamp 1681685098
transform 1 0 1020 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1681685098
transform 1 0 1044 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1278
timestamp 1681685098
transform 1 0 956 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_894
timestamp 1681685098
transform 1 0 964 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1681685098
transform 1 0 996 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1279
timestamp 1681685098
transform 1 0 1044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1681685098
transform 1 0 964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1681685098
transform 1 0 996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1681685098
transform 1 0 1060 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_906
timestamp 1681685098
transform 1 0 1148 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1347
timestamp 1681685098
transform 1 0 1148 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_876
timestamp 1681685098
transform 1 0 1180 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_1262
timestamp 1681685098
transform 1 0 1196 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1681685098
transform 1 0 1164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1681685098
transform 1 0 1188 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1681685098
transform 1 0 1164 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_907
timestamp 1681685098
transform 1 0 1196 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1282
timestamp 1681685098
transform 1 0 1236 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_896
timestamp 1681685098
transform 1 0 1252 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1320
timestamp 1681685098
transform 1 0 1252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1681685098
transform 1 0 1268 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_882
timestamp 1681685098
transform 1 0 1388 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1263
timestamp 1681685098
transform 1 0 1316 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_897
timestamp 1681685098
transform 1 0 1412 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1681685098
transform 1 0 1316 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1681685098
transform 1 0 1428 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_1322
timestamp 1681685098
transform 1 0 1404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1681685098
transform 1 0 1412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1681685098
transform 1 0 1420 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_883
timestamp 1681685098
transform 1 0 1532 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1283
timestamp 1681685098
transform 1 0 1444 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_898
timestamp 1681685098
transform 1 0 1492 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1284
timestamp 1681685098
transform 1 0 1532 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_909
timestamp 1681685098
transform 1 0 1468 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1325
timestamp 1681685098
transform 1 0 1492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1681685098
transform 1 0 1532 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_918
timestamp 1681685098
transform 1 0 1492 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_1285
timestamp 1681685098
transform 1 0 1556 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_899
timestamp 1681685098
transform 1 0 1580 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_1286
timestamp 1681685098
transform 1 0 1588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1681685098
transform 1 0 1596 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_919
timestamp 1681685098
transform 1 0 1596 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_1348
timestamp 1681685098
transform 1 0 1612 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_933
timestamp 1681685098
transform 1 0 1612 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1287
timestamp 1681685098
transform 1 0 1628 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_910
timestamp 1681685098
transform 1 0 1636 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1328
timestamp 1681685098
transform 1 0 1652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1681685098
transform 1 0 1668 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_911
timestamp 1681685098
transform 1 0 1676 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1288
timestamp 1681685098
transform 1 0 1692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1681685098
transform 1 0 1684 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_920
timestamp 1681685098
transform 1 0 1652 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1681685098
transform 1 0 1684 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1681685098
transform 1 0 1668 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1681685098
transform 1 0 1716 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1289
timestamp 1681685098
transform 1 0 1716 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_935
timestamp 1681685098
transform 1 0 1716 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1331
timestamp 1681685098
transform 1 0 1780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1681685098
transform 1 0 1788 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_945
timestamp 1681685098
transform 1 0 1780 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_1349
timestamp 1681685098
transform 1 0 1812 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1681685098
transform 1 0 1828 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_936
timestamp 1681685098
transform 1 0 1820 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1290
timestamp 1681685098
transform 1 0 1860 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_922
timestamp 1681685098
transform 1 0 1852 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1681685098
transform 1 0 1876 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_1351
timestamp 1681685098
transform 1 0 1876 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_884
timestamp 1681685098
transform 1 0 1916 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1291
timestamp 1681685098
transform 1 0 1916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1681685098
transform 1 0 1900 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1681685098
transform 1 0 1908 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_923
timestamp 1681685098
transform 1 0 1908 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_1335
timestamp 1681685098
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_893
timestamp 1681685098
transform 1 0 1964 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_1292
timestamp 1681685098
transform 1 0 1956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1681685098
transform 1 0 1956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1681685098
transform 1 0 1964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1681685098
transform 1 0 1972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1681685098
transform 1 0 1948 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_937
timestamp 1681685098
transform 1 0 1948 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1681685098
transform 1 0 1980 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1681685098
transform 1 0 1972 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1353
timestamp 1681685098
transform 1 0 1980 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_885
timestamp 1681685098
transform 1 0 1996 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_1354
timestamp 1681685098
transform 1 0 2004 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_946
timestamp 1681685098
transform 1 0 2004 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_1293
timestamp 1681685098
transform 1 0 2020 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1681685098
transform 1 0 2028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1681685098
transform 1 0 2036 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1681685098
transform 1 0 2052 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_924
timestamp 1681685098
transform 1 0 2028 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_1295
timestamp 1681685098
transform 1 0 2060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1681685098
transform 1 0 2068 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_939
timestamp 1681685098
transform 1 0 2068 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_1341
timestamp 1681685098
transform 1 0 2084 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1681685098
transform 1 0 2100 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_925
timestamp 1681685098
transform 1 0 2084 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_1356
timestamp 1681685098
transform 1 0 2092 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_940
timestamp 1681685098
transform 1 0 2100 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1681685098
transform 1 0 2092 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_1296
timestamp 1681685098
transform 1 0 2116 0 1 535
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_30
timestamp 1681685098
transform 1 0 24 0 1 470
box -10 -3 10 3
use FILL  FILL_1301
timestamp 1681685098
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1681685098
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1681685098
transform 1 0 88 0 -1 570
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1681685098
transform 1 0 96 0 -1 570
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1681685098
transform 1 0 104 0 -1 570
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1681685098
transform 1 0 112 0 -1 570
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1681685098
transform 1 0 120 0 -1 570
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1681685098
transform 1 0 128 0 -1 570
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1681685098
transform 1 0 136 0 -1 570
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1681685098
transform 1 0 144 0 -1 570
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1681685098
transform 1 0 152 0 -1 570
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1681685098
transform 1 0 160 0 -1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_17
timestamp 1681685098
transform 1 0 168 0 -1 570
box -8 -3 64 105
use FILL  FILL_1325
timestamp 1681685098
transform 1 0 224 0 -1 570
box -8 -3 16 105
use AND2X2  AND2X2_28
timestamp 1681685098
transform 1 0 232 0 -1 570
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1681685098
transform -1 0 360 0 -1 570
box -8 -3 104 105
use OAI21X1  OAI21X1_58
timestamp 1681685098
transform -1 0 392 0 -1 570
box -8 -3 34 105
use AOI22X1  AOI22X1_8
timestamp 1681685098
transform -1 0 432 0 -1 570
box -8 -3 46 105
use FILL  FILL_1326
timestamp 1681685098
transform 1 0 432 0 -1 570
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1681685098
transform 1 0 440 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1681685098
transform 1 0 448 0 -1 570
box -8 -3 104 105
use OR2X1  OR2X1_40
timestamp 1681685098
transform -1 0 576 0 -1 570
box -8 -3 40 105
use XNOR2X1  XNOR2X1_38
timestamp 1681685098
transform 1 0 576 0 -1 570
box -8 -3 64 105
use FILL  FILL_1338
timestamp 1681685098
transform 1 0 632 0 -1 570
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1681685098
transform 1 0 640 0 -1 570
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1681685098
transform 1 0 648 0 -1 570
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1681685098
transform 1 0 656 0 -1 570
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1681685098
transform 1 0 664 0 -1 570
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1681685098
transform 1 0 672 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_46
timestamp 1681685098
transform 1 0 680 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1681685098
transform 1 0 704 0 -1 570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1681685098
transform -1 0 824 0 -1 570
box -8 -3 104 105
use FILL  FILL_1361
timestamp 1681685098
transform 1 0 824 0 -1 570
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1681685098
transform 1 0 832 0 -1 570
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1681685098
transform 1 0 840 0 -1 570
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1681685098
transform 1 0 848 0 -1 570
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1681685098
transform 1 0 856 0 -1 570
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1681685098
transform 1 0 864 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_47
timestamp 1681685098
transform -1 0 896 0 -1 570
box -8 -3 32 105
use FILL  FILL_1374
timestamp 1681685098
transform 1 0 896 0 -1 570
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1681685098
transform 1 0 904 0 -1 570
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1681685098
transform 1 0 912 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_60
timestamp 1681685098
transform 1 0 920 0 -1 570
box -8 -3 34 105
use FILL  FILL_1392
timestamp 1681685098
transform 1 0 952 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1681685098
transform -1 0 1056 0 -1 570
box -8 -3 104 105
use FILL  FILL_1393
timestamp 1681685098
transform 1 0 1056 0 -1 570
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1681685098
transform 1 0 1064 0 -1 570
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1681685098
transform 1 0 1072 0 -1 570
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1681685098
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1681685098
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1681685098
transform 1 0 1096 0 -1 570
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1681685098
transform 1 0 1104 0 -1 570
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1681685098
transform 1 0 1112 0 -1 570
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1681685098
transform 1 0 1120 0 -1 570
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1681685098
transform 1 0 1128 0 -1 570
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1681685098
transform 1 0 1136 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_49
timestamp 1681685098
transform -1 0 1168 0 -1 570
box -8 -3 32 105
use OR2X1  OR2X1_41
timestamp 1681685098
transform -1 0 1200 0 -1 570
box -8 -3 40 105
use FILL  FILL_1416
timestamp 1681685098
transform 1 0 1200 0 -1 570
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1681685098
transform 1 0 1208 0 -1 570
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1681685098
transform 1 0 1216 0 -1 570
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1681685098
transform 1 0 1224 0 -1 570
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1681685098
transform 1 0 1232 0 -1 570
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1681685098
transform 1 0 1240 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_64
timestamp 1681685098
transform 1 0 1248 0 -1 570
box -9 -3 26 105
use FILL  FILL_1428
timestamp 1681685098
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1681685098
transform 1 0 1272 0 -1 570
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1681685098
transform 1 0 1280 0 -1 570
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1681685098
transform 1 0 1288 0 -1 570
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1681685098
transform 1 0 1296 0 -1 570
box -8 -3 16 105
use FAX1  FAX1_6
timestamp 1681685098
transform -1 0 1424 0 -1 570
box -5 -3 126 105
use FILL  FILL_1450
timestamp 1681685098
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1681685098
transform 1 0 1432 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_65
timestamp 1681685098
transform 1 0 1528 0 -1 570
box -9 -3 26 105
use FILL  FILL_1451
timestamp 1681685098
transform 1 0 1544 0 -1 570
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1681685098
transform 1 0 1552 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_61
timestamp 1681685098
transform 1 0 1560 0 -1 570
box -8 -3 34 105
use FILL  FILL_1459
timestamp 1681685098
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1681685098
transform 1 0 1600 0 -1 570
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1681685098
transform 1 0 1608 0 -1 570
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1681685098
transform 1 0 1616 0 -1 570
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1681685098
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1681685098
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1681685098
transform 1 0 1640 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_9
timestamp 1681685098
transform 1 0 1648 0 -1 570
box -8 -3 46 105
use FILL  FILL_1475
timestamp 1681685098
transform 1 0 1688 0 -1 570
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1681685098
transform 1 0 1696 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_66
timestamp 1681685098
transform -1 0 1720 0 -1 570
box -9 -3 26 105
use FILL  FILL_1481
timestamp 1681685098
transform 1 0 1720 0 -1 570
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1681685098
transform 1 0 1728 0 -1 570
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1681685098
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1681685098
transform 1 0 1744 0 -1 570
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1681685098
transform 1 0 1752 0 -1 570
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1681685098
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1681685098
transform 1 0 1768 0 -1 570
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1681685098
transform 1 0 1776 0 -1 570
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1681685098
transform 1 0 1784 0 -1 570
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1681685098
transform 1 0 1792 0 -1 570
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1681685098
transform 1 0 1800 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_52
timestamp 1681685098
transform -1 0 1832 0 -1 570
box -8 -3 32 105
use FILL  FILL_1502
timestamp 1681685098
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1681685098
transform 1 0 1840 0 -1 570
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1681685098
transform 1 0 1848 0 -1 570
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1681685098
transform 1 0 1856 0 -1 570
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1681685098
transform 1 0 1864 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_53
timestamp 1681685098
transform -1 0 1896 0 -1 570
box -8 -3 32 105
use FILL  FILL_1507
timestamp 1681685098
transform 1 0 1896 0 -1 570
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1681685098
transform 1 0 1904 0 -1 570
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1681685098
transform 1 0 1912 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_62
timestamp 1681685098
transform 1 0 1920 0 -1 570
box -8 -3 34 105
use INVX2  INVX2_68
timestamp 1681685098
transform 1 0 1952 0 -1 570
box -9 -3 26 105
use FILL  FILL_1514
timestamp 1681685098
transform 1 0 1968 0 -1 570
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1681685098
transform 1 0 1976 0 -1 570
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1681685098
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1681685098
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_948
timestamp 1681685098
transform 1 0 2020 0 1 475
box -3 -3 3 3
use NAND2X1  NAND2X1_54
timestamp 1681685098
transform -1 0 2024 0 -1 570
box -8 -3 32 105
use M3_M2  M3_M2_949
timestamp 1681685098
transform 1 0 2060 0 1 475
box -3 -3 3 3
use OAI21X1  OAI21X1_63
timestamp 1681685098
transform 1 0 2024 0 -1 570
box -8 -3 34 105
use FILL  FILL_1518
timestamp 1681685098
transform 1 0 2056 0 -1 570
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1681685098
transform 1 0 2064 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_69
timestamp 1681685098
transform 1 0 2072 0 -1 570
box -9 -3 26 105
use NAND2X1  NAND2X1_55
timestamp 1681685098
transform -1 0 2112 0 -1 570
box -8 -3 32 105
use FILL  FILL_1520
timestamp 1681685098
transform 1 0 2112 0 -1 570
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1681685098
transform 1 0 2120 0 -1 570
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1681685098
transform 1 0 2128 0 -1 570
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1681685098
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_31
timestamp 1681685098
transform 1 0 2194 0 1 470
box -10 -3 10 3
use M2_M1  M2_M1_1394
timestamp 1681685098
transform 1 0 84 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1681685098
transform 1 0 148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1681685098
transform 1 0 132 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1681685098
transform 1 0 140 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_980
timestamp 1681685098
transform 1 0 140 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1681685098
transform 1 0 156 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1370
timestamp 1681685098
transform 1 0 164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1681685098
transform 1 0 180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1681685098
transform 1 0 188 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_981
timestamp 1681685098
transform 1 0 188 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1681685098
transform 1 0 236 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1398
timestamp 1681685098
transform 1 0 236 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_950
timestamp 1681685098
transform 1 0 260 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1681685098
transform 1 0 324 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1681685098
transform 1 0 364 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1681685098
transform 1 0 388 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1357
timestamp 1681685098
transform 1 0 372 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1681685098
transform 1 0 260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1681685098
transform 1 0 268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1681685098
transform 1 0 324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1681685098
transform 1 0 348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1681685098
transform 1 0 364 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_960
timestamp 1681685098
transform 1 0 380 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1681685098
transform 1 0 404 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1681685098
transform 1 0 372 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1401
timestamp 1681685098
transform 1 0 396 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_970
timestamp 1681685098
transform 1 0 404 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1402
timestamp 1681685098
transform 1 0 412 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_983
timestamp 1681685098
transform 1 0 396 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1403
timestamp 1681685098
transform 1 0 484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1681685098
transform 1 0 492 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_971
timestamp 1681685098
transform 1 0 508 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1404
timestamp 1681685098
transform 1 0 516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1681685098
transform 1 0 532 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_984
timestamp 1681685098
transform 1 0 532 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1375
timestamp 1681685098
transform 1 0 580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1681685098
transform 1 0 604 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1681685098
transform 1 0 628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1681685098
transform 1 0 620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1681685098
transform 1 0 636 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_985
timestamp 1681685098
transform 1 0 636 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1408
timestamp 1681685098
transform 1 0 684 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_993
timestamp 1681685098
transform 1 0 676 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1681685098
transform 1 0 708 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1409
timestamp 1681685098
transform 1 0 732 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_962
timestamp 1681685098
transform 1 0 788 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1410
timestamp 1681685098
transform 1 0 780 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_972
timestamp 1681685098
transform 1 0 844 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1411
timestamp 1681685098
transform 1 0 852 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_963
timestamp 1681685098
transform 1 0 876 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1412
timestamp 1681685098
transform 1 0 876 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1681685098
transform 1 0 908 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_973
timestamp 1681685098
transform 1 0 916 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1377
timestamp 1681685098
transform 1 0 932 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_994
timestamp 1681685098
transform 1 0 948 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1413
timestamp 1681685098
transform 1 0 964 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1681685098
transform 1 0 980 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1681685098
transform 1 0 1020 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_964
timestamp 1681685098
transform 1 0 1044 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1415
timestamp 1681685098
transform 1 0 1068 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_987
timestamp 1681685098
transform 1 0 1068 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1681685098
transform 1 0 1044 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1681685098
transform 1 0 1108 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1416
timestamp 1681685098
transform 1 0 1116 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_965
timestamp 1681685098
transform 1 0 1140 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1360
timestamp 1681685098
transform 1 0 1172 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1681685098
transform 1 0 1148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1681685098
transform 1 0 1156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1681685098
transform 1 0 1172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1681685098
transform 1 0 1172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1681685098
transform 1 0 1220 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1681685098
transform 1 0 1252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1681685098
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_975
timestamp 1681685098
transform 1 0 1300 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1418
timestamp 1681685098
transform 1 0 1364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1681685098
transform 1 0 1356 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_988
timestamp 1681685098
transform 1 0 1364 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1681685098
transform 1 0 1356 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1384
timestamp 1681685098
transform 1 0 1428 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_966
timestamp 1681685098
transform 1 0 1436 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1419
timestamp 1681685098
transform 1 0 1420 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1681685098
transform 1 0 1428 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1681685098
transform 1 0 1452 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_952
timestamp 1681685098
transform 1 0 1476 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1361
timestamp 1681685098
transform 1 0 1476 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1681685098
transform 1 0 1468 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1681685098
transform 1 0 1492 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_953
timestamp 1681685098
transform 1 0 1516 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_1386
timestamp 1681685098
transform 1 0 1516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1681685098
transform 1 0 1508 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_976
timestamp 1681685098
transform 1 0 1516 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1681685098
transform 1 0 1556 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1424
timestamp 1681685098
transform 1 0 1524 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1681685098
transform 1 0 1532 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_989
timestamp 1681685098
transform 1 0 1508 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1426
timestamp 1681685098
transform 1 0 1588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1681685098
transform 1 0 1604 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1681685098
transform 1 0 1652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1681685098
transform 1 0 1700 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1681685098
transform 1 0 1708 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1681685098
transform 1 0 1716 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_968
timestamp 1681685098
transform 1 0 1700 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1428
timestamp 1681685098
transform 1 0 1676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1681685098
transform 1 0 1684 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_977
timestamp 1681685098
transform 1 0 1692 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1681685098
transform 1 0 1684 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1681685098
transform 1 0 1724 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_1388
timestamp 1681685098
transform 1 0 1740 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_978
timestamp 1681685098
transform 1 0 1740 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_1430
timestamp 1681685098
transform 1 0 1756 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_997
timestamp 1681685098
transform 1 0 1756 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1365
timestamp 1681685098
transform 1 0 1788 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1681685098
transform 1 0 1788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1681685098
transform 1 0 1796 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_991
timestamp 1681685098
transform 1 0 1788 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_1389
timestamp 1681685098
transform 1 0 1820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1681685098
transform 1 0 1836 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1681685098
transform 1 0 1844 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_998
timestamp 1681685098
transform 1 0 1836 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1366
timestamp 1681685098
transform 1 0 1876 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_999
timestamp 1681685098
transform 1 0 1860 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1390
timestamp 1681685098
transform 1 0 1900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1681685098
transform 1 0 1884 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1681685098
transform 1 0 1908 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_992
timestamp 1681685098
transform 1 0 1900 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1681685098
transform 1 0 1908 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1681685098
transform 1 0 1956 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1681685098
transform 1 0 2004 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_1367
timestamp 1681685098
transform 1 0 2068 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1681685098
transform 1 0 2004 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1681685098
transform 1 0 2060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1681685098
transform 1 0 1980 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1681685098
transform 1 0 2092 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1681685098
transform 1 0 2100 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_979
timestamp 1681685098
transform 1 0 2092 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1681685098
transform 1 0 2084 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_1438
timestamp 1681685098
transform 1 0 2108 0 1 405
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_32
timestamp 1681685098
transform 1 0 48 0 1 370
box -10 -3 10 3
use FILL  FILL_1524
timestamp 1681685098
transform 1 0 72 0 1 370
box -8 -3 16 105
use XOR2X1  XOR2X1_18
timestamp 1681685098
transform 1 0 80 0 1 370
box -8 -3 64 105
use FILL  FILL_1526
timestamp 1681685098
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1681685098
transform 1 0 144 0 1 370
box -8 -3 16 105
use AND2X2  AND2X2_31
timestamp 1681685098
transform 1 0 152 0 1 370
box -8 -3 40 105
use XOR2X1  XOR2X1_19
timestamp 1681685098
transform 1 0 184 0 1 370
box -8 -3 64 105
use FILL  FILL_1532
timestamp 1681685098
transform 1 0 240 0 1 370
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1681685098
transform 1 0 248 0 1 370
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1681685098
transform 1 0 256 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1681685098
transform -1 0 360 0 1 370
box -8 -3 104 105
use FILL  FILL_1538
timestamp 1681685098
transform 1 0 360 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_64
timestamp 1681685098
transform -1 0 400 0 1 370
box -8 -3 34 105
use INVX2  INVX2_70
timestamp 1681685098
transform -1 0 416 0 1 370
box -9 -3 26 105
use FILL  FILL_1539
timestamp 1681685098
transform 1 0 416 0 1 370
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1681685098
transform 1 0 424 0 1 370
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1681685098
transform 1 0 432 0 1 370
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1681685098
transform 1 0 440 0 1 370
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1681685098
transform 1 0 448 0 1 370
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1681685098
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1681685098
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1681685098
transform 1 0 472 0 1 370
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1681685098
transform 1 0 480 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_65
timestamp 1681685098
transform -1 0 520 0 1 370
box -8 -3 34 105
use INVX2  INVX2_71
timestamp 1681685098
transform -1 0 536 0 1 370
box -9 -3 26 105
use FILL  FILL_1571
timestamp 1681685098
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1681685098
transform 1 0 544 0 1 370
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1681685098
transform 1 0 552 0 1 370
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1681685098
transform 1 0 560 0 1 370
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1681685098
transform 1 0 568 0 1 370
box -8 -3 16 105
use OR2X1  OR2X1_42
timestamp 1681685098
transform -1 0 608 0 1 370
box -8 -3 40 105
use FILL  FILL_1582
timestamp 1681685098
transform 1 0 608 0 1 370
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1681685098
transform 1 0 616 0 1 370
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1681685098
transform 1 0 624 0 1 370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_39
timestamp 1681685098
transform -1 0 688 0 1 370
box -8 -3 64 105
use FILL  FILL_1585
timestamp 1681685098
transform 1 0 688 0 1 370
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1681685098
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1681685098
transform 1 0 704 0 1 370
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1681685098
transform 1 0 712 0 1 370
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1681685098
transform 1 0 720 0 1 370
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1681685098
transform 1 0 728 0 1 370
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1681685098
transform 1 0 736 0 1 370
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1681685098
transform 1 0 744 0 1 370
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1681685098
transform 1 0 752 0 1 370
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1681685098
transform 1 0 760 0 1 370
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1681685098
transform 1 0 768 0 1 370
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1681685098
transform 1 0 776 0 1 370
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1681685098
transform 1 0 784 0 1 370
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1681685098
transform 1 0 792 0 1 370
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1681685098
transform 1 0 800 0 1 370
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1681685098
transform 1 0 808 0 1 370
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1681685098
transform 1 0 816 0 1 370
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1681685098
transform 1 0 824 0 1 370
box -8 -3 16 105
use INVX2  INVX2_72
timestamp 1681685098
transform 1 0 832 0 1 370
box -9 -3 26 105
use OAI21X1  OAI21X1_66
timestamp 1681685098
transform 1 0 848 0 1 370
box -8 -3 34 105
use FILL  FILL_1620
timestamp 1681685098
transform 1 0 880 0 1 370
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1681685098
transform 1 0 888 0 1 370
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1681685098
transform 1 0 896 0 1 370
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1681685098
transform 1 0 904 0 1 370
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1681685098
transform 1 0 912 0 1 370
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1681685098
transform 1 0 920 0 1 370
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1681685098
transform 1 0 928 0 1 370
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1681685098
transform 1 0 936 0 1 370
box -8 -3 16 105
use INVX2  INVX2_73
timestamp 1681685098
transform -1 0 960 0 1 370
box -9 -3 26 105
use FILL  FILL_1636
timestamp 1681685098
transform 1 0 960 0 1 370
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1681685098
transform 1 0 968 0 1 370
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1681685098
transform 1 0 976 0 1 370
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1681685098
transform 1 0 984 0 1 370
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1681685098
transform 1 0 992 0 1 370
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1681685098
transform 1 0 1000 0 1 370
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1681685098
transform 1 0 1008 0 1 370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_42
timestamp 1681685098
transform -1 0 1072 0 1 370
box -8 -3 64 105
use FILL  FILL_1648
timestamp 1681685098
transform 1 0 1072 0 1 370
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1681685098
transform 1 0 1080 0 1 370
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1681685098
transform 1 0 1088 0 1 370
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1681685098
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1681685098
transform 1 0 1104 0 1 370
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1681685098
transform 1 0 1112 0 1 370
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1681685098
transform 1 0 1120 0 1 370
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1681685098
transform 1 0 1128 0 1 370
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1681685098
transform 1 0 1136 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_1002
timestamp 1681685098
transform 1 0 1180 0 1 375
box -3 -3 3 3
use OAI21X1  OAI21X1_67
timestamp 1681685098
transform 1 0 1144 0 1 370
box -8 -3 34 105
use INVX2  INVX2_74
timestamp 1681685098
transform -1 0 1192 0 1 370
box -9 -3 26 105
use FILL  FILL_1667
timestamp 1681685098
transform 1 0 1192 0 1 370
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1681685098
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1681685098
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1681685098
transform 1 0 1216 0 1 370
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1681685098
transform 1 0 1224 0 1 370
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1681685098
transform 1 0 1232 0 1 370
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1681685098
transform 1 0 1240 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_1003
timestamp 1681685098
transform 1 0 1308 0 1 375
box -3 -3 3 3
use FAX1  FAX1_7
timestamp 1681685098
transform 1 0 1248 0 1 370
box -5 -3 126 105
use FILL  FILL_1677
timestamp 1681685098
transform 1 0 1368 0 1 370
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1681685098
transform 1 0 1376 0 1 370
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1681685098
transform 1 0 1384 0 1 370
box -8 -3 16 105
use INVX2  INVX2_75
timestamp 1681685098
transform -1 0 1408 0 1 370
box -9 -3 26 105
use FILL  FILL_1692
timestamp 1681685098
transform 1 0 1408 0 1 370
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1681685098
transform 1 0 1416 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_68
timestamp 1681685098
transform 1 0 1424 0 1 370
box -8 -3 34 105
use FILL  FILL_1694
timestamp 1681685098
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1681685098
transform 1 0 1464 0 1 370
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1681685098
transform 1 0 1472 0 1 370
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1681685098
transform 1 0 1480 0 1 370
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1681685098
transform 1 0 1488 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_13
timestamp 1681685098
transform 1 0 1496 0 1 370
box -8 -3 46 105
use XOR2X1  XOR2X1_21
timestamp 1681685098
transform -1 0 1592 0 1 370
box -8 -3 64 105
use FILL  FILL_1700
timestamp 1681685098
transform 1 0 1592 0 1 370
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1681685098
transform 1 0 1600 0 1 370
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1681685098
transform 1 0 1608 0 1 370
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1681685098
transform 1 0 1616 0 1 370
box -8 -3 16 105
use XOR2X1  XOR2X1_22
timestamp 1681685098
transform -1 0 1680 0 1 370
box -8 -3 64 105
use NAND2X1  NAND2X1_56
timestamp 1681685098
transform 1 0 1680 0 1 370
box -8 -3 32 105
use FILL  FILL_1712
timestamp 1681685098
transform 1 0 1704 0 1 370
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1681685098
transform 1 0 1712 0 1 370
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1681685098
transform 1 0 1720 0 1 370
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1681685098
transform 1 0 1728 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_58
timestamp 1681685098
transform -1 0 1760 0 1 370
box -8 -3 32 105
use FILL  FILL_1727
timestamp 1681685098
transform 1 0 1760 0 1 370
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1681685098
transform 1 0 1768 0 1 370
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1681685098
transform 1 0 1776 0 1 370
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1681685098
transform 1 0 1784 0 1 370
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1681685098
transform 1 0 1792 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_69
timestamp 1681685098
transform -1 0 1832 0 1 370
box -8 -3 34 105
use FILL  FILL_1737
timestamp 1681685098
transform 1 0 1832 0 1 370
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1681685098
transform 1 0 1840 0 1 370
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1681685098
transform 1 0 1848 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_59
timestamp 1681685098
transform 1 0 1856 0 1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_70
timestamp 1681685098
transform -1 0 1912 0 1 370
box -8 -3 34 105
use FILL  FILL_1740
timestamp 1681685098
transform 1 0 1912 0 1 370
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1681685098
transform 1 0 1920 0 1 370
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1681685098
transform 1 0 1928 0 1 370
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1681685098
transform 1 0 1936 0 1 370
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1681685098
transform 1 0 1944 0 1 370
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1681685098
transform 1 0 1952 0 1 370
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1681685098
transform 1 0 1960 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1681685098
transform 1 0 1968 0 1 370
box -8 -3 104 105
use FILL  FILL_1757
timestamp 1681685098
transform 1 0 2064 0 1 370
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1681685098
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1681685098
transform 1 0 2080 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_60
timestamp 1681685098
transform -1 0 2112 0 1 370
box -8 -3 32 105
use FILL  FILL_1760
timestamp 1681685098
transform 1 0 2112 0 1 370
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1681685098
transform 1 0 2120 0 1 370
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1681685098
transform 1 0 2128 0 1 370
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1681685098
transform 1 0 2136 0 1 370
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_33
timestamp 1681685098
transform 1 0 2170 0 1 370
box -10 -3 10 3
use M2_M1  M2_M1_1476
timestamp 1681685098
transform 1 0 84 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1681685098
transform 1 0 124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1681685098
transform 1 0 116 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1040
timestamp 1681685098
transform 1 0 116 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1681685098
transform 1 0 148 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1447
timestamp 1681685098
transform 1 0 148 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1681685098
transform 1 0 172 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1041
timestamp 1681685098
transform 1 0 172 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1681685098
transform 1 0 156 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1681685098
transform 1 0 212 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1681685098
transform 1 0 204 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1448
timestamp 1681685098
transform 1 0 212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1681685098
transform 1 0 204 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1024
timestamp 1681685098
transform 1 0 244 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1480
timestamp 1681685098
transform 1 0 236 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1005
timestamp 1681685098
transform 1 0 268 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_1449
timestamp 1681685098
transform 1 0 260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1681685098
transform 1 0 252 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1042
timestamp 1681685098
transform 1 0 260 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1681685098
transform 1 0 252 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_1450
timestamp 1681685098
transform 1 0 380 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1006
timestamp 1681685098
transform 1 0 412 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1681685098
transform 1 0 412 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_1451
timestamp 1681685098
transform 1 0 412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1681685098
transform 1 0 396 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1050
timestamp 1681685098
transform 1 0 380 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1681685098
transform 1 0 404 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_1483
timestamp 1681685098
transform 1 0 428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1681685098
transform 1 0 444 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1043
timestamp 1681685098
transform 1 0 444 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1681685098
transform 1 0 492 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1485
timestamp 1681685098
transform 1 0 516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1681685098
transform 1 0 540 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1007
timestamp 1681685098
transform 1 0 564 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_1452
timestamp 1681685098
transform 1 0 556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1681685098
transform 1 0 564 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1008
timestamp 1681685098
transform 1 0 604 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1681685098
transform 1 0 612 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_1454
timestamp 1681685098
transform 1 0 620 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1039
timestamp 1681685098
transform 1 0 636 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1442
timestamp 1681685098
transform 1 0 676 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1681685098
transform 1 0 684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1681685098
transform 1 0 780 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1681685098
transform 1 0 812 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_1025
timestamp 1681685098
transform 1 0 820 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1456
timestamp 1681685098
transform 1 0 820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1681685098
transform 1 0 812 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1026
timestamp 1681685098
transform 1 0 876 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1457
timestamp 1681685098
transform 1 0 876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1681685098
transform 1 0 844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1681685098
transform 1 0 980 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_1009
timestamp 1681685098
transform 1 0 1036 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1681685098
transform 1 0 1028 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1458
timestamp 1681685098
transform 1 0 1028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1681685098
transform 1 0 1036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1681685098
transform 1 0 1052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1681685098
transform 1 0 1028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1681685098
transform 1 0 1044 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1044
timestamp 1681685098
transform 1 0 1028 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1681685098
transform 1 0 1068 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1491
timestamp 1681685098
transform 1 0 1084 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1015
timestamp 1681685098
transform 1 0 1116 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1681685098
transform 1 0 1140 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1461
timestamp 1681685098
transform 1 0 1140 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1681685098
transform 1 0 1228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1681685098
transform 1 0 1172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1681685098
transform 1 0 1220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1681685098
transform 1 0 1284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1681685098
transform 1 0 1300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1681685098
transform 1 0 1308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1681685098
transform 1 0 1324 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1045
timestamp 1681685098
transform 1 0 1324 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_1464
timestamp 1681685098
transform 1 0 1356 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1016
timestamp 1681685098
transform 1 0 1428 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1681685098
transform 1 0 1396 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1681685098
transform 1 0 1436 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1465
timestamp 1681685098
transform 1 0 1396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1681685098
transform 1 0 1444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1681685098
transform 1 0 1476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1681685098
transform 1 0 1484 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1046
timestamp 1681685098
transform 1 0 1492 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_1500
timestamp 1681685098
transform 1 0 1516 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1032
timestamp 1681685098
transform 1 0 1564 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1466
timestamp 1681685098
transform 1 0 1564 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_1033
timestamp 1681685098
transform 1 0 1588 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1501
timestamp 1681685098
transform 1 0 1588 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1010
timestamp 1681685098
transform 1 0 1684 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_1467
timestamp 1681685098
transform 1 0 1668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1681685098
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1681685098
transform 1 0 1708 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_1034
timestamp 1681685098
transform 1 0 1772 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1502
timestamp 1681685098
transform 1 0 1772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1681685098
transform 1 0 1788 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1681685098
transform 1 0 1788 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1017
timestamp 1681685098
transform 1 0 1924 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_1470
timestamp 1681685098
transform 1 0 1924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1681685098
transform 1 0 1844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1681685098
transform 1 0 1884 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1011
timestamp 1681685098
transform 1 0 2076 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1681685098
transform 1 0 1980 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1681685098
transform 1 0 1996 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1681685098
transform 1 0 1980 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1681685098
transform 1 0 2044 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1681685098
transform 1 0 2108 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1681685098
transform 1 0 2092 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1681685098
transform 1 0 2116 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_1471
timestamp 1681685098
transform 1 0 1980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1681685098
transform 1 0 1996 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1681685098
transform 1 0 2084 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1681685098
transform 1 0 1972 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1047
timestamp 1681685098
transform 1 0 1972 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1681685098
transform 1 0 2108 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1474
timestamp 1681685098
transform 1 0 2108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1681685098
transform 1 0 2116 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1681685098
transform 1 0 2044 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1681685098
transform 1 0 2076 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1681685098
transform 1 0 2092 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1681685098
transform 1 0 2108 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1681685098
transform 1 0 2132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_1052
timestamp 1681685098
transform 1 0 2132 0 1 305
box -3 -3 3 3
use top_module_VIA0  top_module_VIA0_34
timestamp 1681685098
transform 1 0 24 0 1 270
box -10 -3 10 3
use FILL  FILL_1525
timestamp 1681685098
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1681685098
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1681685098
transform 1 0 88 0 -1 370
box -8 -3 16 105
use AND2X2  AND2X2_30
timestamp 1681685098
transform -1 0 128 0 -1 370
box -8 -3 40 105
use FILL  FILL_1529
timestamp 1681685098
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1681685098
transform 1 0 136 0 -1 370
box -8 -3 16 105
use XOR2X1  XOR2X1_20
timestamp 1681685098
transform 1 0 144 0 -1 370
box -8 -3 64 105
use FILL  FILL_1534
timestamp 1681685098
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1681685098
transform 1 0 208 0 -1 370
box -8 -3 16 105
use AND2X2  AND2X2_32
timestamp 1681685098
transform -1 0 248 0 -1 370
box -8 -3 40 105
use FILL  FILL_1536
timestamp 1681685098
transform 1 0 248 0 -1 370
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1681685098
transform 1 0 256 0 -1 370
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1681685098
transform 1 0 264 0 -1 370
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1681685098
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1681685098
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1681685098
transform 1 0 288 0 -1 370
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1681685098
transform 1 0 296 0 -1 370
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1681685098
transform 1 0 304 0 -1 370
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1681685098
transform 1 0 312 0 -1 370
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1681685098
transform 1 0 320 0 -1 370
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1681685098
transform 1 0 328 0 -1 370
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1681685098
transform 1 0 336 0 -1 370
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1681685098
transform 1 0 344 0 -1 370
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1681685098
transform 1 0 352 0 -1 370
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1681685098
transform 1 0 360 0 -1 370
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1681685098
transform 1 0 368 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_10
timestamp 1681685098
transform -1 0 416 0 -1 370
box -8 -3 46 105
use FILL  FILL_1555
timestamp 1681685098
transform 1 0 416 0 -1 370
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1681685098
transform 1 0 424 0 -1 370
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1681685098
transform 1 0 432 0 -1 370
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1681685098
transform 1 0 440 0 -1 370
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1681685098
transform 1 0 448 0 -1 370
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1681685098
transform 1 0 456 0 -1 370
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1681685098
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1681685098
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1681685098
transform 1 0 480 0 -1 370
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1681685098
transform 1 0 488 0 -1 370
box -8 -3 16 105
use AND2X2  AND2X2_33
timestamp 1681685098
transform -1 0 528 0 -1 370
box -8 -3 40 105
use FILL  FILL_1574
timestamp 1681685098
transform 1 0 528 0 -1 370
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1681685098
transform 1 0 536 0 -1 370
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1681685098
transform 1 0 544 0 -1 370
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1681685098
transform 1 0 552 0 -1 370
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1681685098
transform 1 0 560 0 -1 370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_40
timestamp 1681685098
transform -1 0 624 0 -1 370
box -8 -3 64 105
use FILL  FILL_1587
timestamp 1681685098
transform 1 0 624 0 -1 370
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1681685098
transform 1 0 632 0 -1 370
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1681685098
transform 1 0 640 0 -1 370
box -8 -3 16 105
use OR2X1  OR2X1_43
timestamp 1681685098
transform -1 0 680 0 -1 370
box -8 -3 40 105
use FILL  FILL_1590
timestamp 1681685098
transform 1 0 680 0 -1 370
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1681685098
transform 1 0 688 0 -1 370
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1681685098
transform 1 0 696 0 -1 370
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1681685098
transform 1 0 704 0 -1 370
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1681685098
transform 1 0 712 0 -1 370
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1681685098
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1681685098
transform 1 0 728 0 -1 370
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1681685098
transform 1 0 736 0 -1 370
box -8 -3 16 105
use OR2X1  OR2X1_44
timestamp 1681685098
transform -1 0 776 0 -1 370
box -8 -3 40 105
use FILL  FILL_1609
timestamp 1681685098
transform 1 0 776 0 -1 370
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1681685098
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1681685098
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1681685098
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1681685098
transform 1 0 808 0 -1 370
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1681685098
transform 1 0 816 0 -1 370
box -8 -3 16 105
use XNOR2X1  XNOR2X1_41
timestamp 1681685098
transform -1 0 880 0 -1 370
box -8 -3 64 105
use FILL  FILL_1622
timestamp 1681685098
transform 1 0 880 0 -1 370
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1681685098
transform 1 0 888 0 -1 370
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1681685098
transform 1 0 896 0 -1 370
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1681685098
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1681685098
transform 1 0 912 0 -1 370
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1681685098
transform 1 0 920 0 -1 370
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1681685098
transform 1 0 928 0 -1 370
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1681685098
transform 1 0 936 0 -1 370
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1681685098
transform 1 0 944 0 -1 370
box -8 -3 16 105
use OR2X1  OR2X1_45
timestamp 1681685098
transform -1 0 984 0 -1 370
box -8 -3 40 105
use FILL  FILL_1642
timestamp 1681685098
transform 1 0 984 0 -1 370
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1681685098
transform 1 0 992 0 -1 370
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1681685098
transform 1 0 1000 0 -1 370
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1681685098
transform 1 0 1008 0 -1 370
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1681685098
transform 1 0 1016 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_11
timestamp 1681685098
transform 1 0 1024 0 -1 370
box -8 -3 46 105
use FILL  FILL_1651
timestamp 1681685098
transform 1 0 1064 0 -1 370
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1681685098
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1681685098
transform 1 0 1080 0 -1 370
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1681685098
transform 1 0 1088 0 -1 370
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1681685098
transform 1 0 1096 0 -1 370
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1681685098
transform 1 0 1104 0 -1 370
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1681685098
transform 1 0 1112 0 -1 370
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1681685098
transform 1 0 1120 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1681685098
transform 1 0 1128 0 -1 370
box -8 -3 104 105
use FILL  FILL_1672
timestamp 1681685098
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1681685098
transform 1 0 1232 0 -1 370
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1681685098
transform 1 0 1240 0 -1 370
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1681685098
transform 1 0 1248 0 -1 370
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1681685098
transform 1 0 1256 0 -1 370
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1681685098
transform 1 0 1264 0 -1 370
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1681685098
transform 1 0 1272 0 -1 370
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1681685098
transform 1 0 1280 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_12
timestamp 1681685098
transform -1 0 1328 0 -1 370
box -8 -3 46 105
use FILL  FILL_1683
timestamp 1681685098
transform 1 0 1328 0 -1 370
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1681685098
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1681685098
transform 1 0 1344 0 -1 370
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1681685098
transform 1 0 1352 0 -1 370
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1681685098
transform 1 0 1360 0 -1 370
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1681685098
transform 1 0 1368 0 -1 370
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1681685098
transform 1 0 1376 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1681685098
transform 1 0 1384 0 -1 370
box -8 -3 104 105
use FILL  FILL_1698
timestamp 1681685098
transform 1 0 1480 0 -1 370
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1681685098
transform 1 0 1488 0 -1 370
box -8 -3 16 105
use AND2X2  AND2X2_34
timestamp 1681685098
transform -1 0 1528 0 -1 370
box -8 -3 40 105
use FILL  FILL_1703
timestamp 1681685098
transform 1 0 1528 0 -1 370
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1681685098
transform 1 0 1536 0 -1 370
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1681685098
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1681685098
transform 1 0 1552 0 -1 370
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1681685098
transform 1 0 1560 0 -1 370
box -8 -3 16 105
use AND2X2  AND2X2_35
timestamp 1681685098
transform -1 0 1600 0 -1 370
box -8 -3 40 105
use FILL  FILL_1708
timestamp 1681685098
transform 1 0 1600 0 -1 370
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1681685098
transform 1 0 1608 0 -1 370
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1681685098
transform 1 0 1616 0 -1 370
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1681685098
transform 1 0 1624 0 -1 370
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1681685098
transform 1 0 1632 0 -1 370
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1681685098
transform 1 0 1640 0 -1 370
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1681685098
transform 1 0 1648 0 -1 370
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1681685098
transform 1 0 1656 0 -1 370
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1681685098
transform 1 0 1664 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_57
timestamp 1681685098
transform 1 0 1672 0 -1 370
box -8 -3 32 105
use FILL  FILL_1720
timestamp 1681685098
transform 1 0 1696 0 -1 370
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1681685098
transform 1 0 1704 0 -1 370
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1681685098
transform 1 0 1712 0 -1 370
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1681685098
transform 1 0 1720 0 -1 370
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1681685098
transform 1 0 1728 0 -1 370
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1681685098
transform 1 0 1736 0 -1 370
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1681685098
transform 1 0 1744 0 -1 370
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1681685098
transform 1 0 1752 0 -1 370
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1681685098
transform 1 0 1760 0 -1 370
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1681685098
transform 1 0 1768 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_76
timestamp 1681685098
transform -1 0 1792 0 -1 370
box -9 -3 26 105
use FILL  FILL_1745
timestamp 1681685098
transform 1 0 1792 0 -1 370
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1681685098
transform 1 0 1800 0 -1 370
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1681685098
transform 1 0 1808 0 -1 370
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1681685098
transform 1 0 1816 0 -1 370
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1681685098
transform 1 0 1824 0 -1 370
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1681685098
transform 1 0 1832 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1681685098
transform -1 0 1936 0 -1 370
box -8 -3 104 105
use FILL  FILL_1751
timestamp 1681685098
transform 1 0 1936 0 -1 370
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1681685098
transform 1 0 1944 0 -1 370
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1681685098
transform 1 0 1952 0 -1 370
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1681685098
transform 1 0 1960 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_77
timestamp 1681685098
transform -1 0 1984 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1681685098
transform 1 0 1984 0 -1 370
box -8 -3 104 105
use OAI21X1  OAI21X1_71
timestamp 1681685098
transform 1 0 2080 0 -1 370
box -8 -3 34 105
use INVX2  INVX2_78
timestamp 1681685098
transform 1 0 2112 0 -1 370
box -9 -3 26 105
use FILL  FILL_1764
timestamp 1681685098
transform 1 0 2128 0 -1 370
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1681685098
transform 1 0 2136 0 -1 370
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_35
timestamp 1681685098
transform 1 0 2194 0 1 270
box -10 -3 10 3
use M3_M2  M3_M2_1067
timestamp 1681685098
transform 1 0 76 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1681685098
transform 1 0 116 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1681685098
transform 1 0 140 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1681685098
transform 1 0 100 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1681685098
transform 1 0 132 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1519
timestamp 1681685098
transform 1 0 100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1681685098
transform 1 0 156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1681685098
transform 1 0 76 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1681685098
transform 1 0 124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1681685098
transform 1 0 132 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1054
timestamp 1681685098
transform 1 0 188 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_1561
timestamp 1681685098
transform 1 0 180 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1105
timestamp 1681685098
transform 1 0 156 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1681685098
transform 1 0 188 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1681685098
transform 1 0 212 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1681685098
transform 1 0 236 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1681685098
transform 1 0 268 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1521
timestamp 1681685098
transform 1 0 204 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1681685098
transform 1 0 212 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1069
timestamp 1681685098
transform 1 0 364 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1513
timestamp 1681685098
transform 1 0 364 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1681685098
transform 1 0 268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1681685098
transform 1 0 324 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1070
timestamp 1681685098
transform 1 0 412 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1681685098
transform 1 0 428 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1524
timestamp 1681685098
transform 1 0 380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1681685098
transform 1 0 388 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1681685098
transform 1 0 396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1681685098
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1681685098
transform 1 0 428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1681685098
transform 1 0 260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1681685098
transform 1 0 348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1681685098
transform 1 0 364 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1096
timestamp 1681685098
transform 1 0 324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1681685098
transform 1 0 364 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1566
timestamp 1681685098
transform 1 0 404 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1098
timestamp 1681685098
transform 1 0 404 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1529
timestamp 1681685098
transform 1 0 476 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1060
timestamp 1681685098
transform 1 0 500 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1681685098
transform 1 0 540 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1681685098
transform 1 0 540 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1681685098
transform 1 0 556 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_1567
timestamp 1681685098
transform 1 0 500 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1681685098
transform 1 0 508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1681685098
transform 1 0 556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1681685098
transform 1 0 572 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1099
timestamp 1681685098
transform 1 0 572 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1530
timestamp 1681685098
transform 1 0 588 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1063
timestamp 1681685098
transform 1 0 660 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1681685098
transform 1 0 652 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1531
timestamp 1681685098
transform 1 0 636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1681685098
transform 1 0 652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1681685098
transform 1 0 660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1681685098
transform 1 0 644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1681685098
transform 1 0 724 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1107
timestamp 1681685098
transform 1 0 724 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_1572
timestamp 1681685098
transform 1 0 764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1681685098
transform 1 0 820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1681685098
transform 1 0 812 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1108
timestamp 1681685098
transform 1 0 812 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1681685098
transform 1 0 844 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_1574
timestamp 1681685098
transform 1 0 844 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1100
timestamp 1681685098
transform 1 0 844 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1681685098
transform 1 0 900 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1681685098
transform 1 0 916 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1681685098
transform 1 0 924 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1536
timestamp 1681685098
transform 1 0 892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1681685098
transform 1 0 908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1681685098
transform 1 0 924 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1681685098
transform 1 0 900 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1681685098
transform 1 0 916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1681685098
transform 1 0 948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1681685098
transform 1 0 980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1681685098
transform 1 0 988 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1083
timestamp 1681685098
transform 1 0 1028 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1681685098
transform 1 0 1052 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_1578
timestamp 1681685098
transform 1 0 1044 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1681685098
transform 1 0 1084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1681685098
transform 1 0 1068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1681685098
transform 1 0 1124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1681685098
transform 1 0 1116 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1109
timestamp 1681685098
transform 1 0 1084 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1681685098
transform 1 0 1116 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1681685098
transform 1 0 1180 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1543
timestamp 1681685098
transform 1 0 1180 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1057
timestamp 1681685098
transform 1 0 1228 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1681685098
transform 1 0 1220 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1544
timestamp 1681685098
transform 1 0 1236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1681685098
transform 1 0 1244 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1111
timestamp 1681685098
transform 1 0 1236 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1681685098
transform 1 0 1276 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1545
timestamp 1681685098
transform 1 0 1268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1681685098
transform 1 0 1284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1681685098
transform 1 0 1276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1681685098
transform 1 0 1284 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1087
timestamp 1681685098
transform 1 0 1332 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1547
timestamp 1681685098
transform 1 0 1332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1681685098
transform 1 0 1340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1681685098
transform 1 0 1388 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1089
timestamp 1681685098
transform 1 0 1396 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1681685098
transform 1 0 1420 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1584
timestamp 1681685098
transform 1 0 1428 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1088
timestamp 1681685098
transform 1 0 1484 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1681685098
transform 1 0 1476 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1550
timestamp 1681685098
transform 1 0 1508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1681685098
transform 1 0 1476 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1681685098
transform 1 0 1484 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1681685098
transform 1 0 1532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1681685098
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1681685098
transform 1 0 1564 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1059
timestamp 1681685098
transform 1 0 1620 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_1589
timestamp 1681685098
transform 1 0 1612 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1681685098
transform 1 0 1620 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1066
timestamp 1681685098
transform 1 0 1668 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_1514
timestamp 1681685098
transform 1 0 1700 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1681685098
transform 1 0 1708 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_1094
timestamp 1681685098
transform 1 0 1716 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1553
timestamp 1681685098
transform 1 0 1732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1681685098
transform 1 0 1724 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1101
timestamp 1681685098
transform 1 0 1764 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1592
timestamp 1681685098
transform 1 0 1780 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1071
timestamp 1681685098
transform 1 0 1804 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1515
timestamp 1681685098
transform 1 0 1804 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1681685098
transform 1 0 1836 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1681685098
transform 1 0 1812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1681685098
transform 1 0 1820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1681685098
transform 1 0 1812 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1095
timestamp 1681685098
transform 1 0 1820 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1681685098
transform 1 0 1844 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1556
timestamp 1681685098
transform 1 0 1852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1681685098
transform 1 0 1836 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1112
timestamp 1681685098
transform 1 0 1812 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_1595
timestamp 1681685098
transform 1 0 1860 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1102
timestamp 1681685098
transform 1 0 1852 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1681685098
transform 1 0 1860 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1681685098
transform 1 0 1876 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1681685098
transform 1 0 1908 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1681685098
transform 1 0 1972 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1517
timestamp 1681685098
transform 1 0 1972 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1681685098
transform 1 0 1980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1681685098
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1681685098
transform 1 0 1956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1681685098
transform 1 0 1972 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_1104
timestamp 1681685098
transform 1 0 1956 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1681685098
transform 1 0 1972 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1681685098
transform 1 0 2068 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1681685098
transform 1 0 2100 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1518
timestamp 1681685098
transform 1 0 2100 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1681685098
transform 1 0 2076 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1681685098
transform 1 0 2084 0 1 205
box -2 -2 2 2
use top_module_VIA0  top_module_VIA0_36
timestamp 1681685098
transform 1 0 48 0 1 170
box -10 -3 10 3
use XOR2X1  XOR2X1_23
timestamp 1681685098
transform -1 0 128 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_24
timestamp 1681685098
transform -1 0 184 0 1 170
box -8 -3 64 105
use FILL  FILL_1767
timestamp 1681685098
transform 1 0 184 0 1 170
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1681685098
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1681685098
transform 1 0 200 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_1115
timestamp 1681685098
transform 1 0 268 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_25
timestamp 1681685098
transform -1 0 264 0 1 170
box -8 -3 64 105
use M3_M2  M3_M2_1116
timestamp 1681685098
transform 1 0 340 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_68
timestamp 1681685098
transform -1 0 360 0 1 170
box -8 -3 104 105
use OAI21X1  OAI21X1_72
timestamp 1681685098
transform -1 0 392 0 1 170
box -8 -3 34 105
use AOI22X1  AOI22X1_14
timestamp 1681685098
transform -1 0 432 0 1 170
box -8 -3 46 105
use FILL  FILL_1770
timestamp 1681685098
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1681685098
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1681685098
transform 1 0 448 0 1 170
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1681685098
transform 1 0 456 0 1 170
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1681685098
transform 1 0 464 0 1 170
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1681685098
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1681685098
transform 1 0 480 0 1 170
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1681685098
transform 1 0 488 0 1 170
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1681685098
transform 1 0 496 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_1117
timestamp 1681685098
transform 1 0 564 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_26
timestamp 1681685098
transform -1 0 560 0 1 170
box -8 -3 64 105
use FILL  FILL_1779
timestamp 1681685098
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1681685098
transform 1 0 568 0 1 170
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1681685098
transform 1 0 576 0 1 170
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1681685098
transform 1 0 584 0 1 170
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1681685098
transform 1 0 592 0 1 170
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1681685098
transform 1 0 600 0 1 170
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1681685098
transform 1 0 608 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_15
timestamp 1681685098
transform -1 0 656 0 1 170
box -8 -3 46 105
use FILL  FILL_1807
timestamp 1681685098
transform 1 0 656 0 1 170
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1681685098
transform 1 0 664 0 1 170
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1681685098
transform 1 0 672 0 1 170
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1681685098
transform 1 0 680 0 1 170
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1681685098
transform 1 0 688 0 1 170
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1681685098
transform 1 0 696 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_1118
timestamp 1681685098
transform 1 0 724 0 1 175
box -3 -3 3 3
use AND2X2  AND2X2_41
timestamp 1681685098
transform -1 0 736 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_1119
timestamp 1681685098
transform 1 0 748 0 1 175
box -3 -3 3 3
use FILL  FILL_1817
timestamp 1681685098
transform 1 0 736 0 1 170
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1681685098
transform 1 0 744 0 1 170
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1681685098
transform 1 0 752 0 1 170
box -8 -3 16 105
use XOR2X1  XOR2X1_31
timestamp 1681685098
transform 1 0 760 0 1 170
box -8 -3 64 105
use FILL  FILL_1820
timestamp 1681685098
transform 1 0 816 0 1 170
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1681685098
transform 1 0 824 0 1 170
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1681685098
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1681685098
transform 1 0 840 0 1 170
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1681685098
transform 1 0 848 0 1 170
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1681685098
transform 1 0 856 0 1 170
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1681685098
transform 1 0 864 0 1 170
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1681685098
transform 1 0 872 0 1 170
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1681685098
transform 1 0 880 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_16
timestamp 1681685098
transform -1 0 928 0 1 170
box -8 -3 46 105
use FILL  FILL_1829
timestamp 1681685098
transform 1 0 928 0 1 170
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1681685098
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1681685098
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1681685098
transform 1 0 952 0 1 170
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1681685098
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1681685098
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1681685098
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1681685098
transform 1 0 984 0 1 170
box -8 -3 16 105
use XOR2X1  XOR2X1_34
timestamp 1681685098
transform -1 0 1048 0 1 170
box -8 -3 64 105
use FILL  FILL_1850
timestamp 1681685098
transform 1 0 1048 0 1 170
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1681685098
transform 1 0 1056 0 1 170
box -8 -3 16 105
use XOR2X1  XOR2X1_35
timestamp 1681685098
transform -1 0 1120 0 1 170
box -8 -3 64 105
use FILL  FILL_1852
timestamp 1681685098
transform 1 0 1120 0 1 170
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1681685098
transform 1 0 1128 0 1 170
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1681685098
transform 1 0 1136 0 1 170
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1681685098
transform 1 0 1144 0 1 170
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1681685098
transform 1 0 1152 0 1 170
box -8 -3 16 105
use AND2X2  AND2X2_47
timestamp 1681685098
transform -1 0 1192 0 1 170
box -8 -3 40 105
use FILL  FILL_1863
timestamp 1681685098
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1681685098
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1681685098
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1681685098
transform 1 0 1216 0 1 170
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1681685098
transform 1 0 1224 0 1 170
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1681685098
transform 1 0 1232 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_1120
timestamp 1681685098
transform 1 0 1252 0 1 175
box -3 -3 3 3
use FILL  FILL_1869
timestamp 1681685098
transform 1 0 1240 0 1 170
box -8 -3 16 105
use AND2X2  AND2X2_48
timestamp 1681685098
transform -1 0 1280 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_1121
timestamp 1681685098
transform 1 0 1340 0 1 175
box -3 -3 3 3
use XOR2X1  XOR2X1_37
timestamp 1681685098
transform -1 0 1336 0 1 170
box -8 -3 64 105
use FILL  FILL_1870
timestamp 1681685098
transform 1 0 1336 0 1 170
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1681685098
transform 1 0 1344 0 1 170
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1681685098
transform 1 0 1352 0 1 170
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1681685098
transform 1 0 1360 0 1 170
box -8 -3 16 105
use AND2X2  AND2X2_49
timestamp 1681685098
transform -1 0 1400 0 1 170
box -8 -3 40 105
use FILL  FILL_1874
timestamp 1681685098
transform 1 0 1400 0 1 170
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1681685098
transform 1 0 1408 0 1 170
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1681685098
transform 1 0 1416 0 1 170
box -8 -3 16 105
use XOR2X1  XOR2X1_38
timestamp 1681685098
transform 1 0 1424 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_39
timestamp 1681685098
transform -1 0 1536 0 1 170
box -8 -3 64 105
use FILL  FILL_1877
timestamp 1681685098
transform 1 0 1536 0 1 170
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1681685098
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1681685098
transform 1 0 1552 0 1 170
box -8 -3 16 105
use XOR2X1  XOR2X1_42
timestamp 1681685098
transform 1 0 1560 0 1 170
box -8 -3 64 105
use FILL  FILL_1894
timestamp 1681685098
transform 1 0 1616 0 1 170
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1681685098
transform 1 0 1624 0 1 170
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1681685098
transform 1 0 1632 0 1 170
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1681685098
transform 1 0 1640 0 1 170
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1681685098
transform 1 0 1648 0 1 170
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1681685098
transform 1 0 1656 0 1 170
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1681685098
transform 1 0 1664 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_61
timestamp 1681685098
transform 1 0 1672 0 1 170
box -8 -3 32 105
use FILL  FILL_1911
timestamp 1681685098
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1681685098
transform 1 0 1704 0 1 170
box -8 -3 16 105
use INVX2  INVX2_80
timestamp 1681685098
transform -1 0 1728 0 1 170
box -9 -3 26 105
use FILL  FILL_1913
timestamp 1681685098
transform 1 0 1728 0 1 170
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1681685098
transform 1 0 1736 0 1 170
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1681685098
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1681685098
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1681685098
transform 1 0 1760 0 1 170
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1681685098
transform 1 0 1768 0 1 170
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1681685098
transform 1 0 1776 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_63
timestamp 1681685098
transform 1 0 1784 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_73
timestamp 1681685098
transform 1 0 1808 0 1 170
box -8 -3 34 105
use FILL  FILL_1928
timestamp 1681685098
transform 1 0 1840 0 1 170
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1681685098
transform 1 0 1848 0 1 170
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1681685098
transform 1 0 1856 0 1 170
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1681685098
transform 1 0 1864 0 1 170
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1681685098
transform 1 0 1872 0 1 170
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1681685098
transform 1 0 1880 0 1 170
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1681685098
transform 1 0 1888 0 1 170
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1681685098
transform 1 0 1896 0 1 170
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1681685098
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1681685098
transform 1 0 1912 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_74
timestamp 1681685098
transform 1 0 1920 0 1 170
box -8 -3 34 105
use NAND2X1  NAND2X1_64
timestamp 1681685098
transform 1 0 1952 0 1 170
box -8 -3 32 105
use FILL  FILL_1941
timestamp 1681685098
transform 1 0 1976 0 1 170
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1681685098
transform 1 0 1984 0 1 170
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1681685098
transform 1 0 1992 0 1 170
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1681685098
transform 1 0 2000 0 1 170
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1681685098
transform 1 0 2008 0 1 170
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1681685098
transform 1 0 2016 0 1 170
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1681685098
transform 1 0 2024 0 1 170
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1681685098
transform 1 0 2032 0 1 170
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1681685098
transform 1 0 2040 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_75
timestamp 1681685098
transform 1 0 2048 0 1 170
box -8 -3 34 105
use NAND2X1  NAND2X1_65
timestamp 1681685098
transform 1 0 2080 0 1 170
box -8 -3 32 105
use FILL  FILL_1955
timestamp 1681685098
transform 1 0 2104 0 1 170
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1681685098
transform 1 0 2112 0 1 170
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1681685098
transform 1 0 2120 0 1 170
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1681685098
transform 1 0 2128 0 1 170
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1681685098
transform 1 0 2136 0 1 170
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_37
timestamp 1681685098
transform 1 0 2170 0 1 170
box -10 -3 10 3
use top_module_VIA0  top_module_VIA0_38
timestamp 1681685098
transform 1 0 24 0 1 70
box -10 -3 10 3
use FILL  FILL_1781
timestamp 1681685098
transform 1 0 72 0 -1 170
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1681685098
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1681685098
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1681685098
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1681685098
transform 1 0 104 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1129
timestamp 1681685098
transform 1 0 124 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1681685098
transform 1 0 124 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1602
timestamp 1681685098
transform 1 0 124 0 1 135
box -2 -2 2 2
use FILL  FILL_1786
timestamp 1681685098
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1681685098
transform 1 0 120 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1130
timestamp 1681685098
transform 1 0 164 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1639
timestamp 1681685098
transform 1 0 140 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1681685098
transform 1 0 156 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1681685098
transform 1 0 164 0 1 125
box -2 -2 2 2
use AND2X2  AND2X2_36
timestamp 1681685098
transform 1 0 128 0 -1 170
box -8 -3 40 105
use FILL  FILL_1788
timestamp 1681685098
transform 1 0 160 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1147
timestamp 1681685098
transform 1 0 180 0 1 145
box -3 -3 3 3
use FILL  FILL_1789
timestamp 1681685098
transform 1 0 168 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1131
timestamp 1681685098
transform 1 0 204 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1603
timestamp 1681685098
transform 1 0 204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1681685098
transform 1 0 212 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1681685098
transform 1 0 196 0 1 125
box -2 -2 2 2
use AND2X2  AND2X2_37
timestamp 1681685098
transform -1 0 208 0 -1 170
box -8 -3 40 105
use FILL  FILL_1790
timestamp 1681685098
transform 1 0 208 0 -1 170
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1681685098
transform 1 0 216 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1132
timestamp 1681685098
transform 1 0 276 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1681685098
transform 1 0 284 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1605
timestamp 1681685098
transform 1 0 276 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1681685098
transform 1 0 252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1681685098
transform 1 0 284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1681685098
transform 1 0 300 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1170
timestamp 1681685098
transform 1 0 252 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1681685098
transform 1 0 300 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1681685098
transform 1 0 276 0 1 105
box -3 -3 3 3
use XOR2X1  XOR2X1_27
timestamp 1681685098
transform -1 0 280 0 -1 170
box -8 -3 64 105
use AND2X2  AND2X2_38
timestamp 1681685098
transform -1 0 312 0 -1 170
box -8 -3 40 105
use FILL  FILL_1792
timestamp 1681685098
transform 1 0 312 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1149
timestamp 1681685098
transform 1 0 332 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1681685098
transform 1 0 348 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1681685098
transform 1 0 380 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1606
timestamp 1681685098
transform 1 0 332 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1681685098
transform 1 0 340 0 1 135
box -2 -2 2 2
use FILL  FILL_1793
timestamp 1681685098
transform 1 0 320 0 -1 170
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1681685098
transform 1 0 328 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1150
timestamp 1681685098
transform 1 0 404 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1608
timestamp 1681685098
transform 1 0 404 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1681685098
transform 1 0 348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1681685098
transform 1 0 356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1681685098
transform 1 0 380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1681685098
transform 1 0 404 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1172
timestamp 1681685098
transform 1 0 356 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1681685098
transform 1 0 380 0 1 115
box -3 -3 3 3
use INVX2  INVX2_79
timestamp 1681685098
transform 1 0 336 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_1174
timestamp 1681685098
transform 1 0 412 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1681685098
transform 1 0 404 0 1 105
box -3 -3 3 3
use XOR2X1  XOR2X1_28
timestamp 1681685098
transform -1 0 408 0 -1 170
box -8 -3 64 105
use FILL  FILL_1795
timestamp 1681685098
transform 1 0 408 0 -1 170
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1681685098
transform 1 0 416 0 -1 170
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1681685098
transform 1 0 424 0 -1 170
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1681685098
transform 1 0 432 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1151
timestamp 1681685098
transform 1 0 468 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1609
timestamp 1681685098
transform 1 0 468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1681685098
transform 1 0 476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1681685098
transform 1 0 460 0 1 125
box -2 -2 2 2
use AND2X2  AND2X2_39
timestamp 1681685098
transform -1 0 472 0 -1 170
box -8 -3 40 105
use FILL  FILL_1799
timestamp 1681685098
transform 1 0 472 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1152
timestamp 1681685098
transform 1 0 532 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1611
timestamp 1681685098
transform 1 0 532 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1163
timestamp 1681685098
transform 1 0 540 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_1651
timestamp 1681685098
transform 1 0 508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1681685098
transform 1 0 540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1681685098
transform 1 0 556 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1175
timestamp 1681685098
transform 1 0 508 0 1 115
box -3 -3 3 3
use XOR2X1  XOR2X1_29
timestamp 1681685098
transform -1 0 536 0 -1 170
box -8 -3 64 105
use M3_M2  M3_M2_1176
timestamp 1681685098
transform 1 0 556 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1681685098
transform 1 0 572 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1612
timestamp 1681685098
transform 1 0 572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1681685098
transform 1 0 580 0 1 135
box -2 -2 2 2
use AND2X2  AND2X2_40
timestamp 1681685098
transform -1 0 568 0 -1 170
box -8 -3 40 105
use M2_M1  M2_M1_1654
timestamp 1681685098
transform 1 0 588 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1177
timestamp 1681685098
transform 1 0 580 0 1 115
box -3 -3 3 3
use FILL  FILL_1800
timestamp 1681685098
transform 1 0 568 0 -1 170
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1681685098
transform 1 0 576 0 -1 170
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1681685098
transform 1 0 584 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1136
timestamp 1681685098
transform 1 0 644 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1614
timestamp 1681685098
transform 1 0 644 0 1 135
box -2 -2 2 2
use XOR2X1  XOR2X1_30
timestamp 1681685098
transform -1 0 648 0 -1 170
box -8 -3 64 105
use FILL  FILL_1809
timestamp 1681685098
transform 1 0 648 0 -1 170
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1681685098
transform 1 0 656 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1153
timestamp 1681685098
transform 1 0 676 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1655
timestamp 1681685098
transform 1 0 676 0 1 125
box -2 -2 2 2
use FILL  FILL_1812
timestamp 1681685098
transform 1 0 664 0 -1 170
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1681685098
transform 1 0 672 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1656
timestamp 1681685098
transform 1 0 700 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1192
timestamp 1681685098
transform 1 0 700 0 1 105
box -3 -3 3 3
use AND2X2  AND2X2_42
timestamp 1681685098
transform -1 0 712 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_1178
timestamp 1681685098
transform 1 0 724 0 1 115
box -3 -3 3 3
use FILL  FILL_1835
timestamp 1681685098
transform 1 0 712 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1122
timestamp 1681685098
transform 1 0 764 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_1615
timestamp 1681685098
transform 1 0 740 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1166
timestamp 1681685098
transform 1 0 740 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1681685098
transform 1 0 732 0 1 95
box -3 -3 3 3
use FILL  FILL_1836
timestamp 1681685098
transform 1 0 720 0 -1 170
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1681685098
transform 1 0 728 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1154
timestamp 1681685098
transform 1 0 788 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1616
timestamp 1681685098
transform 1 0 788 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_1179
timestamp 1681685098
transform 1 0 756 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1681685098
transform 1 0 804 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1681685098
transform 1 0 828 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1681685098
transform 1 0 820 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1617
timestamp 1681685098
transform 1 0 828 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1681685098
transform 1 0 836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1681685098
transform 1 0 796 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1681685098
transform 1 0 804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1681685098
transform 1 0 820 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1180
timestamp 1681685098
transform 1 0 796 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1681685098
transform 1 0 788 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1681685098
transform 1 0 788 0 1 95
box -3 -3 3 3
use XOR2X1  XOR2X1_32
timestamp 1681685098
transform 1 0 736 0 -1 170
box -8 -3 64 105
use FILL  FILL_1838
timestamp 1681685098
transform 1 0 792 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1139
timestamp 1681685098
transform 1 0 884 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1681685098
transform 1 0 884 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1619
timestamp 1681685098
transform 1 0 884 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1681685098
transform 1 0 860 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1181
timestamp 1681685098
transform 1 0 820 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1681685098
transform 1 0 836 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1681685098
transform 1 0 860 0 1 115
box -3 -3 3 3
use AND2X2  AND2X2_43
timestamp 1681685098
transform -1 0 832 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_1123
timestamp 1681685098
transform 1 0 900 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_1661
timestamp 1681685098
transform 1 0 900 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1184
timestamp 1681685098
transform 1 0 892 0 1 115
box -3 -3 3 3
use XOR2X1  XOR2X1_33
timestamp 1681685098
transform -1 0 888 0 -1 170
box -8 -3 64 105
use FILL  FILL_1839
timestamp 1681685098
transform 1 0 888 0 -1 170
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1681685098
transform 1 0 896 0 -1 170
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1681685098
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1681685098
transform 1 0 912 0 -1 170
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1681685098
transform 1 0 920 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1662
timestamp 1681685098
transform 1 0 948 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1167
timestamp 1681685098
transform 1 0 956 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1663
timestamp 1681685098
transform 1 0 964 0 1 125
box -2 -2 2 2
use AND2X2  AND2X2_44
timestamp 1681685098
transform -1 0 960 0 -1 170
box -8 -3 40 105
use FILL  FILL_1844
timestamp 1681685098
transform 1 0 960 0 -1 170
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1681685098
transform 1 0 968 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1164
timestamp 1681685098
transform 1 0 988 0 1 135
box -3 -3 3 3
use FILL  FILL_1848
timestamp 1681685098
transform 1 0 976 0 -1 170
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1681685098
transform 1 0 984 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1124
timestamp 1681685098
transform 1 0 1004 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_1620
timestamp 1681685098
transform 1 0 1004 0 1 135
box -2 -2 2 2
use FILL  FILL_1857
timestamp 1681685098
transform 1 0 992 0 -1 170
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1681685098
transform 1 0 1000 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1165
timestamp 1681685098
transform 1 0 1028 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_1664
timestamp 1681685098
transform 1 0 1028 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1125
timestamp 1681685098
transform 1 0 1044 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1681685098
transform 1 0 1052 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1681685098
transform 1 0 1044 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1621
timestamp 1681685098
transform 1 0 1052 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1681685098
transform 1 0 1044 0 1 125
box -2 -2 2 2
use AND2X2  AND2X2_45
timestamp 1681685098
transform -1 0 1040 0 -1 170
box -8 -3 40 105
use FILL  FILL_1859
timestamp 1681685098
transform 1 0 1040 0 -1 170
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1681685098
transform 1 0 1048 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1126
timestamp 1681685098
transform 1 0 1124 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1681685098
transform 1 0 1092 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1622
timestamp 1681685098
transform 1 0 1084 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1681685098
transform 1 0 1092 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1681685098
transform 1 0 1076 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1681685098
transform 1 0 1092 0 1 125
box -2 -2 2 2
use AND2X2  AND2X2_46
timestamp 1681685098
transform -1 0 1088 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_1141
timestamp 1681685098
transform 1 0 1140 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1624
timestamp 1681685098
transform 1 0 1140 0 1 135
box -2 -2 2 2
use XOR2X1  XOR2X1_36
timestamp 1681685098
transform -1 0 1144 0 -1 170
box -8 -3 64 105
use FILL  FILL_1861
timestamp 1681685098
transform 1 0 1144 0 -1 170
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1681685098
transform 1 0 1152 0 -1 170
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1681685098
transform 1 0 1160 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1625
timestamp 1681685098
transform 1 0 1180 0 1 135
box -2 -2 2 2
use FILL  FILL_1882
timestamp 1681685098
transform 1 0 1168 0 -1 170
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1681685098
transform 1 0 1176 0 -1 170
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1681685098
transform 1 0 1184 0 -1 170
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1681685098
transform 1 0 1192 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1142
timestamp 1681685098
transform 1 0 1260 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1601
timestamp 1681685098
transform 1 0 1268 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1681685098
transform 1 0 1252 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1681685098
transform 1 0 1260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1681685098
transform 1 0 1228 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1194
timestamp 1681685098
transform 1 0 1228 0 1 105
box -3 -3 3 3
use XOR2X1  XOR2X1_40
timestamp 1681685098
transform -1 0 1256 0 -1 170
box -8 -3 64 105
use M2_M1  M2_M1_1628
timestamp 1681685098
transform 1 0 1372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1681685098
transform 1 0 1356 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1185
timestamp 1681685098
transform 1 0 1356 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1681685098
transform 1 0 1372 0 1 105
box -3 -3 3 3
use FAX1  FAX1_8
timestamp 1681685098
transform -1 0 1376 0 -1 170
box -5 -3 126 105
use FILL  FILL_1886
timestamp 1681685098
transform 1 0 1376 0 -1 170
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1681685098
transform 1 0 1384 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1629
timestamp 1681685098
transform 1 0 1404 0 1 135
box -2 -2 2 2
use FILL  FILL_1888
timestamp 1681685098
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1670
timestamp 1681685098
transform 1 0 1412 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1168
timestamp 1681685098
transform 1 0 1420 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1671
timestamp 1681685098
transform 1 0 1428 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1681685098
transform 1 0 1436 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1196
timestamp 1681685098
transform 1 0 1412 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1681685098
transform 1 0 1436 0 1 115
box -3 -3 3 3
use AND2X2  AND2X2_50
timestamp 1681685098
transform 1 0 1400 0 -1 170
box -8 -3 40 105
use FILL  FILL_1889
timestamp 1681685098
transform 1 0 1432 0 -1 170
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1681685098
transform 1 0 1440 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1143
timestamp 1681685098
transform 1 0 1476 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1630
timestamp 1681685098
transform 1 0 1476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1681685098
transform 1 0 1484 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1681685098
transform 1 0 1468 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1169
timestamp 1681685098
transform 1 0 1484 0 1 125
box -3 -3 3 3
use AND2X2  AND2X2_51
timestamp 1681685098
transform -1 0 1480 0 -1 170
box -8 -3 40 105
use FILL  FILL_1891
timestamp 1681685098
transform 1 0 1480 0 -1 170
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1681685098
transform 1 0 1488 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1144
timestamp 1681685098
transform 1 0 1532 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1632
timestamp 1681685098
transform 1 0 1548 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1681685098
transform 1 0 1564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1681685098
transform 1 0 1548 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1681685098
transform 1 0 1556 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1187
timestamp 1681685098
transform 1 0 1548 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1681685098
transform 1 0 1556 0 1 105
box -3 -3 3 3
use XOR2X1  XOR2X1_41
timestamp 1681685098
transform 1 0 1496 0 -1 170
box -8 -3 64 105
use FILL  FILL_1893
timestamp 1681685098
transform 1 0 1552 0 -1 170
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1681685098
transform 1 0 1560 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1145
timestamp 1681685098
transform 1 0 1596 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1676
timestamp 1681685098
transform 1 0 1580 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1681685098
transform 1 0 1596 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1188
timestamp 1681685098
transform 1 0 1580 0 1 115
box -3 -3 3 3
use AND2X2  AND2X2_52
timestamp 1681685098
transform 1 0 1568 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_1189
timestamp 1681685098
transform 1 0 1612 0 1 115
box -3 -3 3 3
use FILL  FILL_1896
timestamp 1681685098
transform 1 0 1600 0 -1 170
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1681685098
transform 1 0 1608 0 -1 170
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1681685098
transform 1 0 1616 0 -1 170
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1681685098
transform 1 0 1624 0 -1 170
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1681685098
transform 1 0 1632 0 -1 170
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1681685098
transform 1 0 1640 0 -1 170
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1681685098
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1634
timestamp 1681685098
transform 1 0 1668 0 1 135
box -2 -2 2 2
use FILL  FILL_1908
timestamp 1681685098
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1681685098
transform 1 0 1664 0 -1 170
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1681685098
transform 1 0 1672 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1685
timestamp 1681685098
transform 1 0 1700 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_62
timestamp 1681685098
transform 1 0 1680 0 -1 170
box -8 -3 32 105
use FILL  FILL_1915
timestamp 1681685098
transform 1 0 1704 0 -1 170
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1681685098
transform 1 0 1712 0 -1 170
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1681685098
transform 1 0 1720 0 -1 170
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1681685098
transform 1 0 1728 0 -1 170
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1681685098
transform 1 0 1736 0 -1 170
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1681685098
transform 1 0 1744 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1635
timestamp 1681685098
transform 1 0 1764 0 1 135
box -2 -2 2 2
use FILL  FILL_1924
timestamp 1681685098
transform 1 0 1752 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1159
timestamp 1681685098
transform 1 0 1860 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1636
timestamp 1681685098
transform 1 0 1860 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1681685098
transform 1 0 1772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1681685098
transform 1 0 1780 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1681685098
transform 1 0 1836 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1200
timestamp 1681685098
transform 1 0 1780 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1681685098
transform 1 0 1804 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1681685098
transform 1 0 1852 0 1 85
box -3 -3 3 3
use INVX2  INVX2_81
timestamp 1681685098
transform 1 0 1760 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_1203
timestamp 1681685098
transform 1 0 1876 0 1 85
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_69
timestamp 1681685098
transform -1 0 1872 0 -1 170
box -8 -3 104 105
use FILL  FILL_1933
timestamp 1681685098
transform 1 0 1872 0 -1 170
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1681685098
transform 1 0 1880 0 -1 170
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1681685098
transform 1 0 1888 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1160
timestamp 1681685098
transform 1 0 1924 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1681685098
transform 1 0 1988 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1637
timestamp 1681685098
transform 1 0 1988 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1681685098
transform 1 0 1908 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1681685098
transform 1 0 1948 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_1204
timestamp 1681685098
transform 1 0 1908 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1681685098
transform 1 0 1932 0 1 85
box -3 -3 3 3
use FILL  FILL_1945
timestamp 1681685098
transform 1 0 1896 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1681685098
transform -1 0 2000 0 -1 170
box -8 -3 104 105
use FILL  FILL_1946
timestamp 1681685098
transform 1 0 2000 0 -1 170
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1681685098
transform 1 0 2008 0 -1 170
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1681685098
transform 1 0 2016 0 -1 170
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1681685098
transform 1 0 2024 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_1127
timestamp 1681685098
transform 1 0 2084 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1681685098
transform 1 0 2124 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1681685098
transform 1 0 2044 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1638
timestamp 1681685098
transform 1 0 2044 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1681685098
transform 1 0 2076 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1681685098
transform 1 0 2124 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_71
timestamp 1681685098
transform 1 0 2032 0 -1 170
box -8 -3 104 105
use FILL  FILL_1959
timestamp 1681685098
transform 1 0 2128 0 -1 170
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1681685098
transform 1 0 2136 0 -1 170
box -8 -3 16 105
use top_module_VIA0  top_module_VIA0_39
timestamp 1681685098
transform 1 0 2194 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1681685098
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_5
timestamp 1681685098
transform 1 0 2170 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_6
timestamp 1681685098
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_7
timestamp 1681685098
transform 1 0 2194 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal3 2218 1125 2218 1125 4 in_clka
rlabel metal3 2218 865 2218 865 4 in_clkb
rlabel metal3 2218 1075 2218 1075 4 in_restart
rlabel metal2 1420 1 1420 1 4 in_inserted_5
rlabel metal2 1572 1 1572 1 4 in_inserted_1
rlabel metal3 2218 935 2218 935 4 in_inserted_05
rlabel metal3 2218 915 2218 915 4 in_inserted_025
rlabel metal2 1052 2038 1052 2038 4 in_sel_a
rlabel metal2 1036 2038 1036 2038 4 in_sel_b
rlabel metal2 1260 2038 1260 2038 4 in_sel_c
rlabel metal2 1348 2038 1348 2038 4 in_sel_d
rlabel metal3 2218 955 2218 955 4 in_next
rlabel metal3 2218 975 2218 975 4 in_finish
rlabel metal3 2 1125 2 1125 4 out_change[15]
rlabel metal3 2 925 2 925 4 out_change[14]
rlabel metal2 756 1 756 1 4 out_change[13]
rlabel metal2 788 1 788 1 4 out_change[12]
rlabel metal2 676 1 676 1 4 out_change[11]
rlabel metal3 2218 525 2218 525 4 out_change[10]
rlabel metal2 1716 1 1716 1 4 out_change[9]
rlabel metal3 2218 505 2218 505 4 out_change[8]
rlabel metal2 1772 1 1772 1 4 out_change[7]
rlabel metal3 2218 325 2218 325 4 out_change[6]
rlabel metal2 1788 1 1788 1 4 out_change[5]
rlabel metal3 2218 305 2218 305 4 out_change[4]
rlabel metal3 2218 545 2218 545 4 out_change[3]
rlabel metal3 2218 615 2218 615 4 out_change[2]
rlabel metal3 2218 725 2218 725 4 out_change[1]
rlabel metal3 2 815 2 815 4 out_change[0]
rlabel metal3 2 1265 2 1265 4 out_stock_a
rlabel metal2 732 2038 732 2038 4 out_stock_b
rlabel metal2 1284 2038 1284 2038 4 out_stock_c
rlabel metal3 2218 1425 2218 1425 4 out_stock_d
rlabel metal2 1140 2038 1140 2038 4 out_csel_a
rlabel metal2 1068 2038 1068 2038 4 out_csel_b
rlabel metal2 1300 2038 1300 2038 4 out_csel_c
rlabel metal2 1436 2038 1436 2038 4 out_csel_d
rlabel metal3 2218 575 2218 575 4 out_change_1[7]
rlabel metal2 1804 1 1804 1 4 out_change_1[6]
rlabel metal3 2218 595 2218 595 4 out_change_1[5]
rlabel metal2 1932 1 1932 1 4 out_change_1[4]
rlabel metal3 2218 165 2218 165 4 out_change_1[3]
rlabel metal2 1852 1 1852 1 4 out_change_1[2]
rlabel metal3 2218 365 2218 365 4 out_change_1[1]
rlabel metal3 2218 475 2218 475 4 out_change_1[0]
rlabel metal3 2218 745 2218 745 4 out_change_05
rlabel metal3 2218 635 2218 635 4 out_change_025
rlabel metal2 1156 2038 1156 2038 4 out_spit_a
rlabel metal2 1004 2038 1004 2038 4 out_spit_b
rlabel metal2 1484 2038 1484 2038 4 out_spit_c
rlabel metal3 2218 1275 2218 1275 4 out_spit_d
rlabel metal3 2218 845 2218 845 4 out_state[1]
rlabel metal3 2218 885 2218 885 4 out_state[0]
rlabel metal1 38 167 38 167 4 gnd
rlabel metal1 14 67 14 67 4 vdd
<< end >>
